
**** 05/08/08 16:20:51 ******* PSpice 15.7.0 (July 2006) ****** ID# 31062456 *

  


 ****     CIRCUIT DESCRIPTION


******************************************************************************







*.subckt mynand3 A B GND Out Vdd



* MAIN CELL: Component pathname : /home/mentor/jack/jaggu
*     
M_MN956 N$14081 N$11345 0 0 n l=2e-06 w=5e-06
M_MN253 N$300 CK N$298 0 n l=2e-06 w=6e-06
M_MN293 N$331 N$327 N$330 0 n l=2e-06 w=6e-06
M_MN292 N$330 CK N$328 0 n l=2e-06 w=6e-06
M_MN291 N$328 N$329 0 0 n l=2e-06 w=6e-06
M_MN344 N$411 N$11347 N$317 0 n l=2e-06 w=5e-06
M_MN13 N$20 N$21 N$23 0 n l=2e-06 w=6e-06
M_MN402 N$11805 N$11794 0 0 n l=2e-06 w=3e-06
M_MN308 N$343 N$340 0 0 n l=2e-06 w=6e-06
M_MN391 N$11570 N$13243 0 0 n l=2e-06 w=5e-06
M_MN390 N$11570 N$13447 N$1674 0 n l=2e-06 w=5e-06
M_MN768 N$11802 N$11796 N$11803 0 n l=2e-06 w=3e-06
M_MN60 0 N$419 N$63 0 n l=2e-06 w=6e-06
M_MN59 N$46 N$421 N$63 0 n l=2e-06 w=6e-06
M_MN58 0 N$417 N$62 0 n l=2e-06 w=6e-06
M_MN57 N$14092 N$420 N$62 0 n l=2e-06 w=6e-06
M_MN70 N$65 N$56 0 0 n l=2e-06 w=5e-06
M_MN69 N$65 N$53 0 0 n l=2e-06 w=5e-06
M_MN71 N$66 N$65 0 0 n l=2e-06 w=5e-06
M_MN77 N$72 N$71 0 0 n l=2e-06 w=5e-06
M_MN76 N$71 N$61 0 0 n l=2e-06 w=5e-06
M_MN75 N$71 N$60 0 0 n l=2e-06 w=5e-06
M_MN80 N$75 N$74 0 0 n l=2e-06 w=5e-06
M_MN79 N$74 N$63 0 0 n l=2e-06 w=5e-06
M_MN78 N$74 N$62 0 0 n l=2e-06 w=5e-06
M_MN951 N$14074 N$11345 0 0 n l=2e-06 w=5e-06
M_MN950 N$14078 N$14074 N$66 0 n l=2e-06 w=5e-06
M_MN949 N$14078 N$11345 0 0 n l=2e-06 w=5e-06
M_MN38 N$43 N$26 0 0 n l=2e-06 w=6e-06
M_MN43 N$3 N$14046 0 0 n l=2e-06 w=6e-06
M_MN42 N$38 N$14092 0 0 n l=2e-06 w=6e-06
M_MN41 N$28 N$14045 0 0 n l=2e-06 w=6e-06
M_MN47 N$13 N$421 N$56 0 n l=2e-06 w=6e-06
M_MN955 N$14080 N$14074 N$72 0 n l=2e-06 w=5e-06
M_MN954 N$14080 N$11345 0 0 n l=2e-06 w=5e-06
M_MN953 N$14079 N$14074 N$415 0 n l=2e-06 w=5e-06
M_MN952 N$14079 N$11345 0 0 n l=2e-06 w=5e-06
M_MN957 N$14081 N$14074 N$75 0 n l=2e-06 w=5e-06
M_MN53 N$14093 N$420 N$60 0 n l=2e-06 w=6e-06
M_MN52 0 N$419 N$59 0 n l=2e-06 w=6e-06
M_MN51 N$36 N$421 N$59 0 n l=2e-06 w=6e-06
M_MN56 0 N$419 N$61 0 n l=2e-06 w=6e-06
M_MN55 N$25 N$421 N$61 0 n l=2e-06 w=6e-06
M_MN22 N$29 N$28 0 0 n l=2e-06 w=6e-06
M_MN28 N$33 N$14 0 0 n l=2e-06 w=6e-06
M_MN27 N$32 N$28 0 0 n l=2e-06 w=6e-06
M_MN26 N$35 N$33 0 0 n l=2e-06 w=6e-06
M_MN25 N$31 N$28 N$35 0 n l=2e-06 w=6e-06
M_MN24 N$34 N$14 0 0 n l=2e-06 w=6e-06
M_MN30 N$17 N$27 0 0 n l=2e-06 w=6e-06
M_MN74 N$415 N$68 0 0 n l=2e-06 w=5e-06
M_MN73 N$68 N$59 0 0 n l=2e-06 w=5e-06
M_MN72 N$68 N$58 0 0 n l=2e-06 w=5e-06
M_MN37 N$42 N$38 0 0 n l=2e-06 w=6e-06
M_MN36 N$45 N$43 0 0 n l=2e-06 w=6e-06
M_MN35 N$41 N$38 N$45 0 n l=2e-06 w=6e-06
M_MN34 N$44 N$26 0 0 n l=2e-06 w=6e-06
M_MN33 N$41 N$42 N$44 0 n l=2e-06 w=6e-06
M_MN40 H_A_Cout N$37 0 0 n l=2e-06 w=6e-06
M_MN39 N$46 N$41 0 0 n l=2e-06 w=6e-06
M_MN364 N$390 N$14096 0 0 n l=2e-06 w=5e-06
M_MN363 N$389 N$409 N$411 0 n l=2e-06 w=5e-06
M_MN362 N$389 N$14096 P4 0 n l=2e-06 w=5e-06
M_MN46 0 N$417 N$53 0 n l=2e-06 w=6e-06
M_MN45 N$14046 N$420 N$53 0 n l=2e-06 w=6e-06
M_MN44 N$16 N$14093 0 0 n l=2e-06 w=6e-06
M_MN50 0 N$417 N$58 0 n l=2e-06 w=6e-06
M_MN49 N$14045 N$420 N$58 0 n l=2e-06 w=6e-06
M_MN48 0 N$419 N$56 0 n l=2e-06 w=6e-06
M_MN54 0 N$417 N$60 0 n l=2e-06 w=6e-06
M_MN20 N$26 N$15 0 0 n l=2e-06 w=6e-06
M_MN19 N$25 N$20 0 0 n l=2e-06 w=6e-06
M_MN23 N$31 N$32 N$34 0 n l=2e-06 w=6e-06
M_MN370 N$395 N$14096 0 0 n l=2e-06 w=5e-06
M_MN7 N$9 N$3 0 0 n l=2e-06 w=6e-06
M_MN357 N$386 N$409 N$372 0 n l=2e-06 w=5e-06
M_MN161 N$182 N$390 0 0 n l=2e-06 w=3e-06
M_MN160 N$181 N$14078 N$182 0 n l=2e-06 w=3e-06
M_MN159 N$180 N$156 0 0 n l=2e-06 w=3e-06
M_MN158 N$180 N$390 0 0 n l=2e-06 w=3e-06
M_MN157 N$180 N$14078 0 0 n l=2e-06 w=3e-06
M_MN29 N$36 N$31 0 0 n l=2e-06 w=6e-06
M_MN32 N$39 N$38 0 0 n l=2e-06 w=6e-06
M_MN31 N$37 N$26 N$39 0 n l=2e-06 w=6e-06
M_MN740 N$11088 N$11327 N$11330 0 n l=2e-06 w=6e-06
M_MN739 N$11330 CK N$11328 0 n l=2e-06 w=6e-06
M_MN738 N$11328 N$11329 0 0 n l=2e-06 w=6e-06
M_MN767 N$11347 N$11345 0 0 n l=2e-06 w=5e-06
M_MN766 N$11345 N$11088 0 0 n l=2e-06 w=5e-06
M_MN747 N$11345 N$11344 0 0 n l=2e-06 w=5e-06
M_MN365 N$390 N$409 N$376 0 n l=2e-06 w=5e-06
M_MN727 N$11322 CK N$11320 0 n l=2e-06 w=6e-06
M_MN726 N$11320 N$11321 N$14096 0 n l=2e-06 w=6e-06
M_MN725 N$11315 CK 0 0 n l=2e-06 w=5e-06
M_MN83 N$81 0 N$85 0 n l=2e-06 w=3e-06
M_MN82 N$85 0 0 0 n l=2e-06 w=3e-06
M_MN81 N$84 N$81 0 0 n l=2e-06 w=3e-06
M_MN271 N$314 CK N$312 0 n l=2e-06 w=6e-06
M_MN270 N$312 N$313 N$250 0 n l=2e-06 w=6e-06
M_MN269 N$306 CK 0 0 n l=2e-06 w=5e-06
M_MN737 N$11329 N$11326 0 0 n l=2e-06 w=6e-06
M_MN310 N$344 CK N$342 0 n l=2e-06 w=6e-06
M_MN309 N$342 N$343 0 0 n l=2e-06 w=6e-06
M_MN350 N$397 N$11347 N$338 0 n l=2e-06 w=5e-06
M_MN349 N$397 N$14095 N$14090 0 n l=2e-06 w=5e-06
M_MN337 N$372 N$14095 N$14084 0 n l=2e-06 w=5e-06
M_MN336 N$14095 N$11347 0 0 n l=2e-06 w=5e-06
M_MN335 N$398 N$11347 N$361 0 n l=2e-06 w=5e-06
M_MN338 N$372 N$11347 N$296 0 n l=2e-06 w=5e-06
M_MN382 N$11779 CK N$11781 0 n l=2e-06 w=6e-06
M_MN387 N$12632 N$11775 0 0 n l=2e-06 w=6e-06
M_MN386 N$12632 N$11780 N$11777 0 n l=2e-06 w=6e-06
M_MN322 N$14086 N$11347 0 0 n l=2e-06 w=5e-06
M_MN321 N$14085 N$348 N$384 0 n l=2e-06 w=5e-06
M_MN320 N$14085 N$11347 0 0 n l=2e-06 w=5e-06
M_MN717 N$11314 N$11315 N$382 0 n l=2e-06 w=6e-06
M_MN186 N$214 N$394 0 0 n l=2e-06 w=3e-06
M_MN185 N$214 N$14080 0 0 n l=2e-06 w=3e-06
M_MN10 N$14 N$2 0 0 n l=2e-06 w=6e-06
M_MN728 N$11323 N$11320 0 0 n l=2e-06 w=6e-06
M_MN327 N$14088 N$11347 0 0 n l=2e-06 w=5e-06
M_MN332 N$14090 N$348 N$338 0 n l=2e-06 w=5e-06
M_MN179 N$207 N$205 0 0 n l=2e-06 w=3e-06
M_MN722 N$14096 N$11315 N$11318 0 n l=2e-06 w=6e-06
M_MN749 N$11334 CK N$11332 0 n l=2e-06 w=6e-06
M_MN378 N$14107 N$11787 0 0 n l=2e-06 w=6e-06
M_MN662 N$1450 N$1485 0 0 n l=2e-06 w=3e-06
M_MN661 N$1435 N$1484 0 0 n l=2e-06 w=3e-06
M_MN693 N$1398 N$1397 0 0 n l=2e-06 w=6e-06
M_MN694 N$1396 CK N$1398 0 n l=2e-06 w=6e-06
M_MN688 N$1401 N$1402 0 0 n l=2e-06 w=6e-06
M_MN702 N$1392 N$1391 0 0 n l=2e-06 w=6e-06
M_MN701 N$1391 N$1394 0 0 n l=2e-06 w=6e-06
M_MN706 N$1389 N$1390 0 0 n l=2e-06 w=6e-06
M_MN705 N$14093 N$1389 0 0 n l=2e-06 w=6e-06
M_MN385 N$11777 CK N$11779 0 n l=2e-06 w=6e-06
M_MN372 N$11784 N$11789 N$11570 0 n l=2e-06 w=6e-06
M_MN176 N$196 N$188 N$197 0 n l=2e-06 w=3e-06
M_MN175 N$199 N$392 0 0 n l=2e-06 w=3e-06
M_MN342 N$374 N$11347 N$310 0 n l=2e-06 w=5e-06
M_MN341 N$374 N$14095 N$14086 0 n l=2e-06 w=5e-06
M_MN188 N$215 N$14080 N$216 0 n l=2e-06 w=3e-06
M_MN187 N$214 N$190 0 0 n l=2e-06 w=3e-06
M_MN110 N$121 0 0 0 n l=2e-06 w=3e-06
M_MN109 N$120 N$118 0 0 n l=2e-06 w=3e-06
M_MN138 N$157 0 0 0 n l=2e-06 w=3e-06
M_MN137 N$156 N$154 0 0 n l=2e-06 w=3e-06
M_MN319 N$14084 N$348 N$296 0 n l=2e-06 w=5e-06
M_MN328 N$14088 N$348 N$324 0 n l=2e-06 w=5e-06
M_MN696 N$14045 N$1395 0 0 n l=2e-06 w=6e-06
M_MN695 N$14045 N$1399 N$1396 0 n l=2e-06 w=6e-06
M_MN659 N$1481 N$1488 0 0 n l=2e-06 w=3e-06
M_MN658 N$1422 N$1426 0 0 n l=2e-06 w=3e-06
M_MN297 N$333 N$334 N$262 0 n l=2e-06 w=6e-06
M_MN333 N$14091 N$348 N$345 0 n l=2e-06 w=5e-06
M_MN12 N$18 N$16 0 0 n l=2e-06 w=6e-06
M_MN11 N$15 N$17 N$18 0 n l=2e-06 w=6e-06
M_MN729 N$11322 N$11323 0 0 n l=2e-06 w=6e-06
M_MN730 N$11324 CK N$11322 0 n l=2e-06 w=6e-06
M_MN672 N$14097 N$1557 N$1467 0 n l=2e-06 w=5e-06
M_MN97 N$100 N$84 N$103 0 n l=2e-06 w=3e-06
M_MN96 N$103 0 0 0 n l=2e-06 w=3e-06
M_MN890 N$14028 N$14040 0 0 n l=2e-06 w=5e-06
M_MN334 N$398 N$14095 OUT8 0 n l=2e-06 w=5e-06
M_MN754 N$382 N$11337 0 0 n l=2e-06 w=6e-06
M_MN724 N$11319 N$11318 0 0 n l=2e-06 w=6e-06
M_MN14 N$23 N$17 0 0 n l=2e-06 w=6e-06
M_MN312 N$345 N$346 0 0 n l=2e-06 w=6e-06
M_MN123 N$138 N$136 0 0 n l=2e-06 w=3e-06
M_MN704 N$14093 N$1393 N$1390 0 n l=2e-06 w=6e-06
M_MN709 N$1386 CK N$1388 0 n l=2e-06 w=6e-06
M_MN296 N$327 CK 0 0 n l=2e-06 w=5e-06
M_MN84 N$86 N$385 0 0 n l=2e-06 w=3e-06
M_MN112 N$122 N$387 0 0 n l=2e-06 w=3e-06
M_MN111 N$118 N$102 N$121 0 n l=2e-06 w=3e-06
M_MN550 N$1529 N$1530 0 0 n l=2e-06 w=5e-06
M_MN549 N$1529 N$14108 N$14107 0 n l=2e-06 w=5e-06
M_MN418 N$1662 N$11809 N$1660 0 n l=2e-06 w=3e-06
M_MN422 N$1651 N$1668 N$1649 0 n l=2e-06 w=3e-06
M_MN421 N$1649 N$11561 0 0 n l=2e-06 w=3e-06
M_MN420 N$1650 N$1651 0 0 n l=2e-06 w=3e-06
M_MN15 N$20 N$16 N$24 0 n l=2e-06 w=6e-06
M_MN697 N$1395 N$1396 0 0 n l=2e-06 w=6e-06
M_MN703 N$1390 CK N$1392 0 n l=2e-06 w=6e-06
M_MN669 N$1504 N$1416 N$1526 0 n l=2e-06 w=5e-06
M_MN674 N$1413 N$1557 0 0 n l=2e-06 w=5e-06
M_MN673 N$14097 N$1413 0 0 n l=2e-06 w=5e-06
M_MN759 N$11341 N$11338 0 0 n l=2e-06 w=6e-06
M_MN758 N$11340 CK N$11338 0 n l=2e-06 w=6e-06
M_MN757 N$11338 N$11339 N$11099 0 n l=2e-06 w=6e-06
M_MN756 N$11333 CK 0 0 n l=2e-06 w=5e-06
M_MN765 N$11339 CK 0 0 n l=2e-06 w=5e-06
M_MN755 N$11337 N$11336 0 0 n l=2e-06 w=6e-06
M_MN770 N$11810 N$11802 0 0 n l=2e-06 w=3e-06
M_MN520 N$1553 N$1558 0 0 n l=2e-06 w=5e-06
M_MN519 N$13857 N$1554 N$1553 0 n l=2e-06 w=5e-06
M_MN723 N$14096 N$11319 0 0 n l=2e-06 w=6e-06
M_MN746 N$11345 N$11099 0 0 n l=2e-06 w=5e-06
M_MN315 OUT8 N$11347 0 0 n l=2e-06 w=5e-06
M_MN347 N$412 N$14095 N$14089 0 n l=2e-06 w=5e-06
M_MN346 N$376 N$11347 N$324 0 n l=2e-06 w=5e-06
M_MN414 N$1661 N$11809 0 0 n l=2e-06 w=3e-06
M_MN413 N$1661 N$1673 0 0 n l=2e-06 w=3e-06
M_MN412 N$1661 N$1654 0 0 n l=2e-06 w=3e-06
M_MN419 N$13038 N$1662 0 0 n l=2e-06 w=3e-06
M_MN389 N$11780 CK 0 0 n l=2e-06 w=5e-06
M_MN479 N$1593 N$13447 N$1654 0 n l=2e-06 w=5e-06
M_MN478 N$11816 N$13243 N$1654 0 n l=2e-06 w=5e-06
M_MN477 N$11816 N$13447 N$11561 0 n l=2e-06 w=5e-06
M_MN518 N$1557 N$11083 0 0 n l=2e-06 w=5e-06
M_MN517 N$1557 N$1558 0 0 n l=2e-06 w=5e-06
M_MN764 N$11343 N$11342 0 0 n l=2e-06 w=6e-06
M_MN763 N$11344 N$11343 0 0 n l=2e-06 w=6e-06
M_MN762 N$11344 N$11339 N$11342 0 n l=2e-06 w=6e-06
M_MN761 N$11342 CK N$11340 0 n l=2e-06 w=6e-06
M_MN760 N$11340 N$11341 0 0 n l=2e-06 w=6e-06
M_MN539 N$14108 N$13857 0 0 n l=2e-06 w=6e-06
M_MN538 N$1544 CK 0 0 n l=2e-06 w=5e-06
M_MN537 N$11083 N$1540 0 0 n l=2e-06 w=6e-06
M_MN558 N$1523 N$1522 N$1521 0 n l=2e-06 w=6e-06
M_MN557 N$1525 N$1530 0 0 n l=2e-06 w=5e-06
M_MN439 N$1634 N$11786 N$1631 0 n l=2e-06 w=3e-06
M_MN438 N$1632 N$1636 0 0 n l=2e-06 w=3e-06
M_MN437 N$1631 N$1636 0 0 n l=2e-06 w=3e-06
M_MN436 N$1634 N$1650 N$1632 0 n l=2e-06 w=3e-06
M_MN470 N$1595 N$13447 N$1599 0 n l=2e-06 w=5e-06
M_MN469 N$13650 N$12835 0 0 n l=2e-06 w=6e-06
M_MN745 N$11345 N$14096 0 0 n l=2e-06 w=5e-06
M_MN744 N$11345 N$382 0 0 n l=2e-06 w=5e-06
M_MN522 N$1549 CK N$1552 0 n l=2e-06 w=6e-06
M_MN417 N$1662 N$1671 N$1661 0 n l=2e-06 w=3e-06
M_MN416 N$1659 N$1673 0 0 n l=2e-06 w=3e-06
M_MN415 N$1660 N$1654 N$1659 0 n l=2e-06 w=3e-06
M_MN499 N$1573 N$1572 N$1595 0 n l=2e-06 w=6e-06
M_MN504 N$12429 N$1572 N$1569 0 n l=2e-06 w=6e-06
M_MN471 N$1595 N$13243 N$11786 0 n l=2e-06 w=5e-06
M_MN476 N$11817 N$13243 N$11561 0 n l=2e-06 w=5e-06
M_MN475 N$11817 N$13447 N$11786 0 n l=2e-06 w=5e-06
M_MN521 N$1552 N$1551 N$13650 0 n l=2e-06 w=6e-06
M_MN487 N$11571 N$1581 0 0 n l=2e-06 w=6e-06
M_MN507 N$1572 CK 0 0 n l=2e-06 w=5e-06
M_MN506 N$12633 N$1569 0 0 n l=2e-06 w=6e-06
M_MN435 N$1632 N$11786 0 0 n l=2e-06 w=3e-06
M_MN523 N$1548 N$1552 0 0 n l=2e-06 w=6e-06
M_MN500 N$1571 CK N$1573 0 n l=2e-06 w=6e-06
M_MN486 N$11571 N$1588 N$1583 0 n l=2e-06 w=6e-06
M_MN483 N$1584 N$1589 0 0 n l=2e-06 w=6e-06
M_MN461 N$13039 N$1611 0 0 n l=2e-06 w=3e-06
M_MN473 N$13650 N$13039 0 0 n l=2e-06 w=5e-06
M_MN432 N$1644 N$1668 N$1642 0 n l=2e-06 w=3e-06
M_MN431 N$1644 N$1651 N$1643 0 n l=2e-06 w=3e-06
M_MN430 N$1641 N$1653 0 0 n l=2e-06 w=3e-06
M_MN429 N$1642 N$11561 N$1641 0 n l=2e-06 w=3e-06
M_MN434 N$1633 N$1634 0 0 n l=2e-06 w=3e-06
M_MN93 N$90 0 N$92 0 n l=2e-06 w=3e-06
M_MN92 N$90 N$81 N$91 0 n l=2e-06 w=3e-06
M_MN91 N$93 N$385 0 0 n l=2e-06 w=3e-06
M_MN90 N$92 0 N$93 0 n l=2e-06 w=3e-06
M_MN89 N$91 0 0 0 n l=2e-06 w=3e-06
M_MN290 N$329 N$326 0 0 n l=2e-06 w=6e-06
M_MN289 N$328 CK N$326 0 n l=2e-06 w=6e-06
M_MN468 N$13650 N$13037 0 0 n l=2e-06 w=6e-06
M_MN467 N$13650 N$13038 0 0 n l=2e-06 w=6e-06
M_MN541 N$1674 N$11813 N$14107 0 n l=2e-06 w=5e-06
M_MN472 N$13243 N$13447 0 0 n l=2e-06 w=5e-06
M_MN445 N$1627 N$1634 N$1626 0 n l=2e-06 w=3e-06
M_MN444 N$1624 N$1636 0 0 n l=2e-06 w=3e-06
M_MN443 N$1625 N$11786 N$1624 0 n l=2e-06 w=3e-06
M_MN388 N$11775 N$11777 0 0 n l=2e-06 w=6e-06
M_MN453 N$9715 N$1599 N$1615 0 n l=2e-06 w=3e-06
M_MN457 N$1609 N$1599 N$1608 0 n l=2e-06 w=3e-06
M_MN456 N$1610 N$1633 0 0 n l=2e-06 w=3e-06
M_MN440 N$1626 N$11786 0 0 n l=2e-06 w=3e-06
M_MN441 N$1626 N$1636 0 0 n l=2e-06 w=3e-06
M_MN442 N$1626 N$1650 0 0 n l=2e-06 w=3e-06
M_MN265 N$309 CK N$307 0 n l=2e-06 w=6e-06
M_MN264 N$307 N$308 0 0 n l=2e-06 w=6e-06
M_MN263 N$308 N$305 0 0 n l=2e-06 w=6e-06
M_MN240 N$417 N$420 0 0 n l=2e-06 w=6e-06
M_MN205 N$230 N$207 N$232 0 n l=2e-06 w=3e-06
M_MN239 N$420 N$279 0 0 n l=2e-06 w=6e-06
M_MN433 N$13037 N$1644 0 0 n l=2e-06 w=3e-06
M_MN590 SK3 N$1497 N$1493 0 n l=2e-06 w=6e-06
M_MN563 SK0 N$1522 N$1517 0 n l=2e-06 w=6e-06
M_MN562 N$1517 CK N$1519 0 n l=2e-06 w=6e-06
M_MN155 N$174 N$390 0 0 n l=2e-06 w=3e-06
M_MN154 N$175 N$390 0 0 n l=2e-06 w=3e-06
M_MN198 N$222 N$14081 N$226 0 n l=2e-06 w=3e-06
M_MN197 N$225 N$395 0 0 n l=2e-06 w=3e-06
M_MN196 N$226 N$395 0 0 n l=2e-06 w=3e-06
M_MN195 N$222 N$207 N$225 0 n l=2e-06 w=3e-06
M_MN194 N$225 N$14081 0 0 n l=2e-06 w=3e-06
M_MN94 N$94 N$90 0 0 n l=2e-06 w=3e-06
M_MN275 N$317 N$313 N$316 0 n l=2e-06 w=6e-06
M_MN274 N$316 CK N$314 0 n l=2e-06 w=6e-06
M_MN273 N$314 N$315 0 0 n l=2e-06 w=6e-06
M_MN246 N$293 N$294 0 0 n l=2e-06 w=6e-06
M_MN298 N$335 CK N$333 0 n l=2e-06 w=6e-06
M_MN86 N$81 0 N$86 0 n l=2e-06 w=3e-06
M_MN85 N$85 N$385 0 0 n l=2e-06 w=3e-06
M_MN113 N$121 N$387 0 0 n l=2e-06 w=3e-06
M_MN142 N$154 0 N$158 0 n l=2e-06 w=3e-06
M_MN141 N$157 N$389 0 0 n l=2e-06 w=3e-06
M_MN409 N$1666 N$1673 0 0 n l=2e-06 w=3e-06
M_MN408 N$1671 N$11809 N$1667 0 n l=2e-06 w=3e-06
M_MN455 N$1610 N$1620 0 0 n l=2e-06 w=3e-06
M_MN454 N$1610 N$1599 0 0 n l=2e-06 w=3e-06
M_MN426 N$1643 N$11561 0 0 n l=2e-06 w=3e-06
M_MN266 N$310 N$306 N$309 0 n l=2e-06 w=6e-06
M_MN492 N$1577 N$1580 0 0 n l=2e-06 w=6e-06
M_MN491 N$1578 CK N$1580 0 n l=2e-06 w=6e-06
M_MN490 N$1580 N$1579 N$11816 0 n l=2e-06 w=6e-06
M_MN489 N$1588 CK 0 0 n l=2e-06 w=5e-06
M_MN261 N$305 N$306 N$246 0 n l=2e-06 w=6e-06
M_MN260 N$299 CK 0 0 n l=2e-06 w=5e-06
M_MN238 N$420 N$386 0 0 n l=2e-06 w=6e-06
M_MN258 N$384 N$304 0 0 n l=2e-06 w=6e-06
M_MN257 N$384 N$299 N$302 0 n l=2e-06 w=6e-06
M_MN282 N$321 N$322 0 0 n l=2e-06 w=6e-06
M_MN281 N$322 N$319 0 0 n l=2e-06 w=6e-06
M_MN532 N$1541 N$1545 0 0 n l=2e-06 w=6e-06
M_MN531 N$1542 CK N$1545 0 n l=2e-06 w=6e-06
M_MN536 N$1554 N$11083 0 0 n l=2e-06 w=6e-06
M_MN503 N$1569 CK N$1571 0 n l=2e-06 w=6e-06
M_MN502 N$1571 N$1570 0 0 n l=2e-06 w=6e-06
M_MN566 N$1522 CK 0 0 n l=2e-06 w=5e-06
M_MN565 N$1515 N$1517 0 0 n l=2e-06 w=6e-06
M_MN564 SK0 N$1515 0 0 n l=2e-06 w=6e-06
M_MN245 N$294 N$291 0 0 n l=2e-06 w=6e-06
M_MN406 N$1668 N$1671 0 0 n l=2e-06 w=3e-06
M_MN244 N$293 CK N$291 0 n l=2e-06 w=6e-06
M_MN243 N$291 N$292 N$237 0 n l=2e-06 w=6e-06
M_MN262 N$307 CK N$305 0 n l=2e-06 w=6e-06
M_MN411 N$1671 N$1654 N$1666 0 n l=2e-06 w=3e-06
M_MN410 N$1667 N$1673 0 0 n l=2e-06 w=3e-06
M_MN576 N$1506 N$1505 N$1504 0 n l=2e-06 w=6e-06
M_MN575 N$1513 CK 0 0 n l=2e-06 w=5e-06
M_MN601 N$1484 N$1557 N$12429 0 n l=2e-06 w=5e-06
M_MN606 N$1475 N$1481 0 0 n l=2e-06 w=3e-06
M_MN605 N$1479 C N$1476 0 n l=2e-06 w=3e-06
M_MN604 N$1476 B0 0 0 n l=2e-06 w=3e-06
M_MN573 SK1 N$1507 0 0 n l=2e-06 w=6e-06
M_MN578 N$1502 N$1506 0 0 n l=2e-06 w=6e-06
M_MN577 N$1503 CK N$1506 0 n l=2e-06 w=6e-06
M_MN581 SK2 N$1505 N$1501 0 n l=2e-06 w=6e-06
M_MN580 N$1501 CK N$1503 0 n l=2e-06 w=6e-06
M_MN495 N$11572 N$1579 N$1576 0 n l=2e-06 w=6e-06
M_MN494 N$1576 CK N$1578 0 n l=2e-06 w=6e-06
M_MN259 N$304 N$302 0 0 n l=2e-06 w=6e-06
M_MN497 N$1574 N$1576 0 0 n l=2e-06 w=6e-06
M_MN496 N$11572 N$1574 0 0 n l=2e-06 w=6e-06
M_MN501 N$1570 N$1573 0 0 n l=2e-06 w=6e-06
M_MN586 N$1495 CK N$1498 0 n l=2e-06 w=6e-06
M_MN622 N$1463 B1 N$1460 0 n l=2e-06 w=3e-06
M_MN589 N$1493 CK N$1495 0 n l=2e-06 w=6e-06
M_MN594 N$1488 N$1557 N$11571 0 n l=2e-06 w=5e-06
M_MN561 N$1519 N$1518 0 0 n l=2e-06 w=6e-06
M_MN592 N$1491 N$1493 0 0 n l=2e-06 w=6e-06
M_MN597 N$1486 N$1557 N$11572 0 n l=2e-06 w=5e-06
M_MN596 N$1489 N$1557 0 0 n l=2e-06 w=5e-06
M_MN569 N$1510 N$1514 0 0 n l=2e-06 w=6e-06
M_MN567 N$1514 N$1513 N$1512 0 n l=2e-06 w=6e-06
M_MN572 SK1 N$1513 N$1509 0 n l=2e-06 w=6e-06
M_MN571 N$1509 CK N$1511 0 n l=2e-06 w=6e-06
M_MN570 N$1511 N$1510 0 0 n l=2e-06 w=6e-06
M_MN602 N$1484 N$1489 0 0 n l=2e-06 w=5e-06
M_MN603 N$1477 N$1479 0 0 n l=2e-06 w=3e-06
M_MN608 N$1479 B0 N$1475 0 n l=2e-06 w=3e-06
M_MN607 N$1476 N$1481 0 0 n l=2e-06 w=3e-06
M_MN611 N$1470 C 0 0 n l=2e-06 w=3e-06
M_MN610 N$1470 N$1481 0 0 n l=2e-06 w=3e-06
M_MN609 N$1470 B0 0 0 n l=2e-06 w=3e-06
M_MN579 N$1503 N$1502 0 0 n l=2e-06 w=6e-06
M_MN585 N$1498 N$1497 N$1496 0 n l=2e-06 w=6e-06
M_MN584 N$1505 CK 0 0 n l=2e-06 w=5e-06
M_MN493 N$1578 N$1577 0 0 n l=2e-06 w=6e-06
M_MN498 N$1579 CK 0 0 n l=2e-06 w=5e-06
M_MN582 SK2 N$1499 0 0 n l=2e-06 w=6e-06
M_MN588 N$1495 N$1494 0 0 n l=2e-06 w=6e-06
M_MN587 N$1494 N$1498 0 0 n l=2e-06 w=6e-06
M_MN649 N$1431 N$1435 0 0 n l=2e-06 w=3e-06
M_MN648 N$1430 N$1435 0 0 n l=2e-06 w=3e-06
M_MN652 N$1425 N$1435 0 0 n l=2e-06 w=3e-06
M_MN651 N$1425 B3 0 0 n l=2e-06 w=3e-06
M_MN621 N$1461 N$1465 0 0 n l=2e-06 w=3e-06
M_MN620 N$1460 N$1465 0 0 n l=2e-06 w=3e-06
M_MN619 N$1463 N$1477 N$1461 0 n l=2e-06 w=3e-06
M_MN593 N$1497 CK 0 0 n l=2e-06 w=5e-06
M_MN629 N$1456 N$1477 N$1454 0 n l=2e-06 w=3e-06
M_MN628 N$1456 N$1463 N$1455 0 n l=2e-06 w=3e-06
M_MN627 N$1453 N$1465 0 0 n l=2e-06 w=3e-06
M_MN595 N$1488 N$1489 0 0 n l=2e-06 w=5e-06
M_MN568 N$1511 CK N$1514 0 n l=2e-06 w=6e-06
M_MN599 N$1485 N$1557 N$12632 0 n l=2e-06 w=5e-06
M_MN598 N$1486 N$1489 0 0 n l=2e-06 w=5e-06
M_MN632 N$1446 B2 0 0 n l=2e-06 w=3e-06
M_MN631 N$1447 N$1448 0 0 n l=2e-06 w=3e-06
M_MN667 N$1512 N$1416 N$1527 0 n l=2e-06 w=5e-06
M_MN666 N$1512 N$1557 N$1486 0 n l=2e-06 w=5e-06
M_MN671 N$1496 N$1416 N$1525 0 n l=2e-06 w=5e-06
M_MN636 N$1448 B2 N$1445 0 n l=2e-06 w=3e-06
M_MN640 N$1439 B2 N$1438 0 n l=2e-06 w=3e-06
M_MN639 N$1440 N$1462 0 0 n l=2e-06 w=3e-06
M_MN638 N$1440 N$1450 0 0 n l=2e-06 w=3e-06
M_MN637 N$1440 B2 0 0 n l=2e-06 w=3e-06
M_MN644 N$1437 N$1441 0 0 n l=2e-06 w=3e-06
M_MN583 N$1499 N$1501 0 0 n l=2e-06 w=6e-06
M_MN615 N$1471 C N$1469 0 n l=2e-06 w=3e-06
M_MN614 N$1471 N$1479 N$1470 0 n l=2e-06 w=3e-06
M_MN613 N$1468 N$1481 0 0 n l=2e-06 w=3e-06
M_MN612 N$1469 B0 N$1468 0 n l=2e-06 w=3e-06
M_MN618 N$1461 B1 0 0 n l=2e-06 w=3e-06
M_MN617 N$1462 N$1463 0 0 n l=2e-06 w=3e-06
M_MN650 N$1433 B3 N$1430 0 n l=2e-06 w=3e-06
M_MN683 N$1403 N$1406 0 0 n l=2e-06 w=6e-06
M_MN682 N$1404 CK N$1406 0 n l=2e-06 w=6e-06
M_MN657 N$1426 N$1447 N$1424 0 n l=2e-06 w=3e-06
M_MN656 N$1426 N$1433 N$1425 0 n l=2e-06 w=3e-06
M_MN655 N$1423 N$1435 0 0 n l=2e-06 w=3e-06
M_MN654 N$1424 B3 N$1423 0 n l=2e-06 w=3e-06
M_MN653 N$1425 N$1447 0 0 n l=2e-06 w=3e-06
M_MN660 N$1465 N$1486 0 0 n l=2e-06 w=3e-06
M_MN626 N$1454 B1 N$1453 0 n l=2e-06 w=3e-06
M_MN625 N$1455 N$1477 0 0 n l=2e-06 w=3e-06
M_MN624 N$1455 N$1465 0 0 n l=2e-06 w=3e-06
M_MN600 N$1485 N$1489 0 0 n l=2e-06 w=5e-06
M_MN630 N$1452 N$1456 0 0 n l=2e-06 w=3e-06
M_MN634 N$1445 N$1450 0 0 n l=2e-06 w=3e-06
M_MN633 N$1448 N$1462 N$1446 0 n l=2e-06 w=3e-06
M_MN668 N$1504 N$1557 N$1485 0 n l=2e-06 w=5e-06
M_MN700 N$1392 CK N$1394 0 n l=2e-06 w=6e-06
M_MN699 N$1394 N$1393 N$1409 0 n l=2e-06 w=6e-06
M_MN698 N$1399 CK 0 0 n l=2e-06 w=5e-06
M_MN670 N$1496 N$1557 N$1484 0 n l=2e-06 w=5e-06
M_MN635 N$1446 N$1450 0 0 n l=2e-06 w=3e-06
M_MN339 N$410 N$14095 N$14085 0 n l=2e-06 w=5e-06
M_MN358 N$387 N$14096 P2 0 n l=2e-06 w=5e-06
M_MN355 N$409 N$14096 0 0 n l=2e-06 w=5e-06
M_MN678 N$1409 N$1413 0 0 n l=2e-06 w=5e-06
M_MN677 N$1409 N$1557 N$1437 0 n l=2e-06 w=5e-06
M_MN616 N$1467 N$1471 0 0 n l=2e-06 w=3e-06
M_MN645 CoutHK_SK N$1433 0 0 n l=2e-06 w=3e-06
M_MN684 N$1404 N$1403 0 0 n l=2e-06 w=6e-06
M_MN715 N$1383 N$1384 0 0 n l=2e-06 w=6e-06
M_MN714 N$14092 N$1383 0 0 n l=2e-06 w=6e-06
M_MN687 N$14046 N$1401 0 0 n l=2e-06 w=6e-06
M_MN397 N$11796 N$1674 N$11798 0 n l=2e-06 w=3e-06
M_MN396 N$11797 N$11794 0 0 n l=2e-06 w=3e-06
M_MN395 N$11798 N$11794 0 0 n l=2e-06 w=3e-06
M_MN394 N$11796 C N$11797 0 n l=2e-06 w=3e-06
M_MN393 N$11797 N$1674 0 0 n l=2e-06 w=3e-06
M_MN235 N$421 N$275 0 0 n l=2e-06 w=6e-06
M_MN234 N$421 N$385 0 0 n l=2e-06 w=6e-06
M_MN623 N$1455 B1 0 0 n l=2e-06 w=3e-06
M_MN665 N$1416 N$1557 0 0 n l=2e-06 w=5e-06
M_MN664 N$1521 N$1416 N$1529 0 n l=2e-06 w=5e-06
M_MN663 N$1521 N$1557 N$1488 0 n l=2e-06 w=5e-06
M_MN555 N$1526 N$1530 0 0 n l=2e-06 w=5e-06
M_MN554 N$1526 N$14108 N$11572 0 n l=2e-06 w=5e-06
M_MN560 N$1518 N$1523 0 0 n l=2e-06 w=6e-06
M_MN559 N$1519 CK N$1523 0 n l=2e-06 w=6e-06
M_MN488 N$1581 N$1583 0 0 n l=2e-06 w=6e-06
M_MN340 N$410 N$11347 N$384 0 n l=2e-06 w=5e-06
M_MN777 OUT0 N$13879 0 0 n l=2e-06 w=3e-06
M_MN776 N$13879 0 N$13881 0 n l=2e-06 w=3e-06
M_MN775 N$13879 N$13870 N$13880 0 n l=2e-06 w=3e-06
M_MN774 N$13882 N$13996 0 0 n l=2e-06 w=3e-06
M_MN574 N$1507 N$1509 0 0 n l=2e-06 w=6e-06
M_MN676 N$1410 N$1413 0 0 n l=2e-06 w=5e-06
M_MN708 N$1388 N$1387 N$1408 0 n l=2e-06 w=6e-06
M_MN707 N$1393 CK 0 0 n l=2e-06 w=5e-06
M_MN713 N$14092 N$1387 N$1384 0 n l=2e-06 w=6e-06
M_MN712 N$1384 CK N$1386 0 n l=2e-06 w=6e-06
M_MN711 N$1386 N$1385 0 0 n l=2e-06 w=6e-06
M_MN511 N$13874 N$13996 0 0 n l=2e-06 w=3e-06
M_MN510 N$13875 N$13996 0 0 n l=2e-06 w=3e-06
M_MN509 N$13870 0 N$13874 0 n l=2e-06 w=3e-06
M_MN508 N$13874 N$14084 0 0 n l=2e-06 w=3e-06
M_MN474 N$13873 N$13870 0 0 n l=2e-06 w=3e-06
M_MN791 OUT1 N$13895 0 0 n l=2e-06 w=3e-06
M_MN790 N$13895 N$13873 N$13897 0 n l=2e-06 w=3e-06
M_MN392 N$11809 N$11796 0 0 n l=2e-06 w=3e-06
M_MN552 N$1527 N$14108 N$11571 0 n l=2e-06 w=5e-06
M_MN551 N$1530 N$14108 0 0 n l=2e-06 w=5e-06
M_MN556 N$1525 N$14108 N$12632 0 n l=2e-06 w=5e-06
M_MN783 N$13887 N$14085 N$13891 0 n l=2e-06 w=3e-06
M_MN782 N$13890 N$14000 0 0 n l=2e-06 w=3e-06
M_MN781 N$13891 N$14000 0 0 n l=2e-06 w=3e-06
M_MN780 N$13887 N$13873 N$13890 0 n l=2e-06 w=3e-06
M_MN779 N$13890 N$14085 0 0 n l=2e-06 w=3e-06
M_MN778 N$13889 N$13887 0 0 n l=2e-06 w=3e-06
M_MN805 OUT2 N$13911 0 0 n l=2e-06 w=3e-06
M_MN516 N$13881 N$14084 N$13882 0 n l=2e-06 w=3e-06
M_MN515 N$13880 0 0 0 n l=2e-06 w=3e-06
M_MN514 N$13880 N$13996 0 0 n l=2e-06 w=3e-06
M_MN553 N$1527 N$1530 0 0 n l=2e-06 w=5e-06
M_MN512 N$13870 N$14084 N$13875 0 n l=2e-06 w=3e-06
M_MN797 N$13903 N$14086 N$13907 0 n l=2e-06 w=3e-06
M_MN796 N$13906 N$14001 0 0 n l=2e-06 w=3e-06
M_MN795 N$13907 N$14001 0 0 n l=2e-06 w=3e-06
M_MN794 N$13903 N$13889 N$13906 0 n l=2e-06 w=3e-06
M_MN793 N$13906 N$14086 0 0 n l=2e-06 w=3e-06
M_MN792 N$13905 N$13903 0 0 n l=2e-06 w=3e-06
M_MN821 N$13938 N$14088 0 0 n l=2e-06 w=3e-06
M_MN820 N$13937 N$13935 0 0 n l=2e-06 w=3e-06
M_MN789 N$13895 N$13887 N$13896 0 n l=2e-06 w=3e-06
M_MN788 N$13898 N$14000 0 0 n l=2e-06 w=3e-06
M_MN787 N$13897 N$14085 N$13898 0 n l=2e-06 w=3e-06
M_MN811 N$13919 N$14087 N$13923 0 n l=2e-06 w=3e-06
M_MN810 N$13922 N$14002 0 0 n l=2e-06 w=3e-06
M_MN809 N$13923 N$14002 0 0 n l=2e-06 w=3e-06
M_MN808 N$13919 N$13905 N$13922 0 n l=2e-06 w=3e-06
M_MN807 N$13922 N$14087 0 0 n l=2e-06 w=3e-06
M_MN806 N$13921 N$13919 0 0 n l=2e-06 w=3e-06
M_MN837 N$13955 N$14004 0 0 n l=2e-06 w=3e-06
M_MN836 N$13951 N$13937 N$13954 0 n l=2e-06 w=3e-06
M_MN835 N$13954 N$14089 0 0 n l=2e-06 w=3e-06
M_MN834 N$13953 N$13951 0 0 n l=2e-06 w=3e-06
M_MN804 N$13911 N$13889 N$13913 0 n l=2e-06 w=3e-06
M_MN803 N$13911 N$13903 N$13912 0 n l=2e-06 w=3e-06
M_MN513 N$13880 N$14084 0 0 n l=2e-06 w=3e-06
M_MN799 N$13912 N$14001 0 0 n l=2e-06 w=3e-06
M_MN798 N$13912 N$14086 0 0 n l=2e-06 w=3e-06
M_MN825 N$13935 N$14088 N$13939 0 n l=2e-06 w=3e-06
M_MN824 N$13938 N$14003 0 0 n l=2e-06 w=3e-06
M_MN823 N$13939 N$14003 0 0 n l=2e-06 w=3e-06
M_MN822 N$13935 N$13921 N$13938 0 n l=2e-06 w=3e-06
M_MN853 N$13967 N$14090 N$13971 0 n l=2e-06 w=3e-06
M_MN852 N$13970 N$14005 0 0 n l=2e-06 w=3e-06
M_MN851 N$13971 N$14005 0 0 n l=2e-06 w=3e-06
M_MN850 N$13967 N$13953 N$13970 0 n l=2e-06 w=3e-06
M_MN849 N$13970 N$14090 0 0 n l=2e-06 w=3e-06
M_MN848 N$13969 N$13967 0 0 n l=2e-06 w=3e-06
M_MN819 OUT3 N$13927 0 0 n l=2e-06 w=3e-06
M_MN786 N$13896 N$13873 0 0 n l=2e-06 w=3e-06
M_MN785 N$13896 N$14000 0 0 n l=2e-06 w=3e-06
M_MN784 N$13896 N$14085 0 0 n l=2e-06 w=3e-06
M_MN815 N$13929 N$14087 N$13930 0 n l=2e-06 w=3e-06
M_MN814 N$13928 N$13905 0 0 n l=2e-06 w=3e-06
M_MN813 N$13928 N$14002 0 0 n l=2e-06 w=3e-06
M_MN812 N$13928 N$14087 0 0 n l=2e-06 w=3e-06
M_MN840 N$13960 N$14089 0 0 n l=2e-06 w=3e-06
M_MN839 N$13951 N$14089 N$13955 0 n l=2e-06 w=3e-06
M_MN838 N$13954 N$14004 0 0 n l=2e-06 w=3e-06
M_MN867 N$13983 N$14091 N$13987 0 n l=2e-06 w=3e-06
M_MN866 N$13986 N$14007 0 0 n l=2e-06 w=3e-06
M_MN865 N$13987 N$14007 0 0 n l=2e-06 w=3e-06
M_MN864 N$13983 N$13969 N$13986 0 n l=2e-06 w=3e-06
M_MN863 N$13986 N$14091 0 0 n l=2e-06 w=3e-06
M_MN862 CARRY_OUT N$13983 0 0 n l=2e-06 w=3e-06
M_MN802 N$13914 N$14001 0 0 n l=2e-06 w=3e-06
M_MN801 N$13913 N$14086 N$13914 0 n l=2e-06 w=3e-06
M_MN800 N$13912 N$13889 0 0 n l=2e-06 w=3e-06
M_MN831 N$13943 N$13935 N$13944 0 n l=2e-06 w=3e-06
M_MN830 N$13946 N$14003 0 0 n l=2e-06 w=3e-06
M_MN829 N$13945 N$14088 N$13946 0 n l=2e-06 w=3e-06
M_MN828 N$13944 N$13921 0 0 n l=2e-06 w=3e-06
M_MN827 N$13944 N$14003 0 0 n l=2e-06 w=3e-06
M_MN826 N$13944 N$14088 0 0 n l=2e-06 w=3e-06
M_MN856 N$13976 N$13953 0 0 n l=2e-06 w=3e-06
M_MN855 N$13976 N$14005 0 0 n l=2e-06 w=3e-06
M_MN854 N$13976 N$14090 0 0 n l=2e-06 w=3e-06
M_MN930 N$14005 N$14006 N$14014 0 n l=2e-06 w=5e-06
M_MN929 N$14006 SK3 0 0 n l=2e-06 w=5e-06
M_MN928 N$14007 SK3 N$14012 0 n l=2e-06 w=5e-06
M_MN933 N$14004 SK3 N$14010 0 n l=2e-06 w=5e-06
M_MN900 N$14021 N$14024 N$14031 0 n l=2e-06 w=5e-06
M_MN899 N$14022 SK1 N$14031 0 n l=2e-06 w=5e-06
M_MN818 N$13927 N$13905 N$13929 0 n l=2e-06 w=3e-06
M_MN817 N$13927 N$13919 N$13928 0 n l=2e-06 w=3e-06
M_MN816 N$13930 N$14002 0 0 n l=2e-06 w=3e-06
M_MN846 N$13959 N$13937 N$13961 0 n l=2e-06 w=3e-06
M_MN845 N$13959 N$13951 N$13960 0 n l=2e-06 w=3e-06
M_MN844 N$13962 N$14004 0 0 n l=2e-06 w=3e-06
M_MN843 N$13961 N$14089 N$13962 0 n l=2e-06 w=3e-06
M_MN842 N$13960 N$13937 0 0 n l=2e-06 w=3e-06
M_MN841 N$13960 N$14004 0 0 n l=2e-06 w=3e-06
M_MN872 N$13994 N$14007 0 0 n l=2e-06 w=3e-06
M_MN871 N$13993 N$14091 N$13994 0 n l=2e-06 w=3e-06
M_MN870 N$13992 N$13969 0 0 n l=2e-06 w=3e-06
M_MN869 N$13992 N$14007 0 0 n l=2e-06 w=3e-06
M_MN868 N$13992 N$14091 0 0 n l=2e-06 w=3e-06
M_MN945 N$14040 N$13857 N$13999 0 n l=2e-06 w=5e-06
M_MN944 N$14040 N$14108 N$11083 0 n l=2e-06 w=5e-06
M_MN948 N$13999 N$13997 0 0 n l=2e-06 w=5e-06
M_MN947 N$13997 N$11347 0 0 n l=2e-06 w=5e-06
M_MN916 N$14013 SK2 N$14020 0 n l=2e-06 w=5e-06
M_MN915 N$14013 N$14015 N$14022 0 n l=2e-06 w=5e-06
M_MN833 OUT4 N$13943 0 0 n l=2e-06 w=3e-06
M_MN832 N$13943 N$13921 N$13945 0 n l=2e-06 w=3e-06
M_MN861 OUT6 N$13975 0 0 n l=2e-06 w=3e-06
M_MN860 N$13975 N$13953 N$13977 0 n l=2e-06 w=3e-06
M_MN859 N$13975 N$13967 N$13976 0 n l=2e-06 w=3e-06
M_MN858 N$13978 N$14005 0 0 n l=2e-06 w=3e-06
M_MN857 N$13977 N$14090 N$13978 0 n l=2e-06 w=3e-06
M_MN922 N$14010 SK2 N$14017 0 n l=2e-06 w=5e-06
M_MN927 N$14007 N$14006 N$14016 0 n l=2e-06 w=5e-06
M_MN926 N$14008 SK2 0 0 n l=2e-06 w=5e-06
M_MN925 N$14008 N$14015 N$14017 0 n l=2e-06 w=5e-06
M_MN222 N$258 N$14095 N$200 0 n l=2e-06 w=5e-06
M_MN299 N$336 N$333 0 0 n l=2e-06 w=6e-06
M_MN231 N$271 N$14095 N$94 0 n l=2e-06 w=5e-06
M_MN905 N$14019 SK1 N$14028 0 n l=2e-06 w=5e-06
M_MN904 N$14019 N$14024 N$14029 0 n l=2e-06 w=5e-06
M_MN903 N$14020 SK1 N$14029 0 n l=2e-06 w=5e-06
M_MN902 N$14020 N$14024 N$14030 0 n l=2e-06 w=5e-06
M_MN908 N$14017 N$14024 N$14027 0 n l=2e-06 w=5e-06
M_MN907 N$14018 SK1 N$14027 0 n l=2e-06 w=5e-06
M_MN938 N$14001 N$14006 N$14010 0 n l=2e-06 w=5e-06
M_MN943 N$13996 SK3 0 0 n l=2e-06 w=5e-06
M_MN942 N$13996 N$14006 N$14008 0 n l=2e-06 w=5e-06
M_MN941 N$14000 SK3 0 0 n l=2e-06 w=5e-06
M_MN946 N$13997 N$11083 0 0 n l=2e-06 w=5e-06
M_MN122 N$130 N$126 0 0 n l=2e-06 w=3e-06
M_MN121 N$126 N$102 N$128 0 n l=2e-06 w=3e-06
M_MN120 N$126 N$118 N$127 0 n l=2e-06 w=3e-06
M_MN119 N$129 N$387 0 0 n l=2e-06 w=3e-06
M_MN118 N$128 0 N$129 0 n l=2e-06 w=3e-06
M_MN88 N$91 N$385 0 0 n l=2e-06 w=3e-06
M_MN87 N$91 0 0 0 n l=2e-06 w=3e-06
M_MN921 N$14010 N$14015 N$14019 0 n l=2e-06 w=5e-06
M_MN920 N$14011 SK2 N$14018 0 n l=2e-06 w=5e-06
M_MN919 N$14011 N$14015 N$14020 0 n l=2e-06 w=5e-06
M_MN918 N$14012 SK2 N$14019 0 n l=2e-06 w=5e-06
M_MN924 N$14009 SK2 0 0 n l=2e-06 w=5e-06
M_MN923 N$14009 N$14015 N$14018 0 n l=2e-06 w=5e-06
M_MN223 N$258 N$265 N$217 0 n l=2e-06 w=5e-06
M_MN210 N$242 N$14095 N$130 0 n l=2e-06 w=5e-06
M_MN170 N$188 N$14079 N$192 0 n l=2e-06 w=3e-06
M_MN108 N$112 N$108 0 0 n l=2e-06 w=3e-06
M_MN107 N$108 N$84 N$110 0 n l=2e-06 w=3e-06
M_MN106 N$108 N$100 N$109 0 n l=2e-06 w=3e-06
M_MN407 N$1667 N$1654 0 0 n l=2e-06 w=3e-06
M_MN206 N$1179 N$230 0 0 n l=2e-06 w=3e-06
M_MN145 N$163 N$138 0 0 n l=2e-06 w=3e-06
M_MN204 N$230 N$222 N$231 0 n l=2e-06 w=3e-06
M_MN203 N$233 N$395 0 0 n l=2e-06 w=3e-06
M_MN202 N$232 N$14081 N$233 0 n l=2e-06 w=3e-06
M_MN201 N$231 N$207 0 0 n l=2e-06 w=3e-06
M_MN200 N$231 N$395 0 0 n l=2e-06 w=3e-06
M_MN237 N$275 N$386 0 0 n l=2e-06 w=6e-06
M_MN236 N$419 N$421 0 0 n l=2e-06 w=6e-06
M_MN288 N$326 N$327 N$258 0 n l=2e-06 w=6e-06
M_MN287 N$320 CK 0 0 n l=2e-06 w=5e-06
M_MN193 Cout N$222 0 0 n l=2e-06 w=3e-06
M_MN184 N$205 N$14080 N$209 0 n l=2e-06 w=3e-06
M_MN183 N$208 N$394 0 0 n l=2e-06 w=3e-06
M_MN182 N$209 N$394 0 0 n l=2e-06 w=3e-06
M_MN181 N$205 N$190 N$208 0 n l=2e-06 w=3e-06
M_MN180 N$208 N$14080 0 0 n l=2e-06 w=3e-06
M_MN95 N$102 N$100 0 0 n l=2e-06 w=3e-06
M_MN692 N$1397 N$1400 0 0 n l=2e-06 w=6e-06
M_MN546 N$11561 N$11813 N$11572 0 n l=2e-06 w=5e-06
M_MN545 N$11561 RST 0 0 n l=2e-06 w=5e-06
M_MN544 N$1654 N$11813 N$11571 0 n l=2e-06 w=5e-06
M_MN543 N$1654 RST 0 0 n l=2e-06 w=5e-06
M_MN542 N$11813 RST 0 0 n l=2e-06 w=5e-06
M_MN377 N$14107 N$11789 N$11790 0 n l=2e-06 w=6e-06
M_MN169 N$191 N$392 0 0 n l=2e-06 w=3e-06
M_MN211 N$242 N$265 N$148 0 n l=2e-06 w=5e-06
M_MN136 N$148 N$144 0 0 n l=2e-06 w=3e-06
M_MN135 N$144 N$120 N$146 0 n l=2e-06 w=3e-06
M_MN134 N$144 N$136 N$145 0 n l=2e-06 w=3e-06
M_MN133 N$147 N$388 0 0 n l=2e-06 w=3e-06
M_MN102 N$109 N$386 0 0 n l=2e-06 w=3e-06
M_MN101 N$109 0 0 0 n l=2e-06 w=3e-06
M_MN105 N$111 N$386 0 0 n l=2e-06 w=3e-06
M_MN104 N$110 0 N$111 0 n l=2e-06 w=3e-06
M_MN103 N$109 N$84 0 0 n l=2e-06 w=3e-06
M_MN330 N$14089 N$348 N$331 0 n l=2e-06 w=5e-06
M_MN307 N$342 CK N$340 0 n l=2e-06 w=6e-06
M_MN306 N$340 N$341 N$266 0 n l=2e-06 w=6e-06
M_MN100 N$100 0 N$104 0 n l=2e-06 w=3e-06
M_MN99 N$103 N$386 0 0 n l=2e-06 w=3e-06
M_MN128 N$136 0 N$140 0 n l=2e-06 w=3e-06
M_MN156 N$171 N$14078 N$175 0 n l=2e-06 w=3e-06
M_MN329 N$14089 N$11347 0 0 n l=2e-06 w=5e-06
M_MN248 N$296 N$292 N$295 0 n l=2e-06 w=6e-06
M_MN247 N$295 CK N$293 0 n l=2e-06 w=6e-06
M_MN217 N$250 N$265 N$183 0 n l=2e-06 w=5e-06
M_MN190 N$213 N$205 N$214 0 n l=2e-06 w=3e-06
M_MN216 N$250 N$14095 N$166 0 n l=2e-06 w=5e-06
M_MN425 N$1651 N$11561 N$1648 0 n l=2e-06 w=3e-06
M_MN424 N$1649 N$1653 0 0 n l=2e-06 w=3e-06
M_MN233 N$265 N$14095 0 0 n l=2e-06 w=5e-06
M_MN189 N$216 N$394 0 0 n l=2e-06 w=3e-06
M_MN208 N$237 N$265 N$130 0 n l=2e-06 w=5e-06
M_MN207 N$237 N$14095 N$112 0 n l=2e-06 w=5e-06
M_MN374 N$11782 N$11784 0 0 n l=2e-06 w=6e-06
M_MN373 N$11783 CK N$11784 0 n l=2e-06 w=6e-06
M_MN63 N$287 N$282 0 0 n l=2e-06 w=6e-06
M_MN64 N$286 N$287 0 0 n l=2e-06 w=6e-06
M_MN65 N$288 CK N$286 0 n l=2e-06 w=6e-06
M_MN191 N$213 N$190 N$215 0 n l=2e-06 w=3e-06
M_MN130 N$145 N$388 0 0 n l=2e-06 w=3e-06
M_MN174 N$198 N$14079 N$199 0 n l=2e-06 w=3e-06
M_MN173 N$197 N$173 0 0 n l=2e-06 w=3e-06
M_MN172 N$197 N$392 0 0 n l=2e-06 w=3e-06
M_MN171 N$197 N$14079 0 0 n l=2e-06 w=3e-06
M_MN214 N$246 N$265 N$166 0 n l=2e-06 w=5e-06
M_MN114 N$118 0 N$122 0 n l=2e-06 w=3e-06
M_MN423 N$1648 N$1653 0 0 n l=2e-06 w=3e-06
M_MN428 N$1643 N$1668 0 0 n l=2e-06 w=3e-06
M_MN427 N$1643 N$1653 0 0 n l=2e-06 w=3e-06
M_MN277 N$318 N$316 0 0 n l=2e-06 w=6e-06
M_MN276 N$317 N$318 0 0 n l=2e-06 w=6e-06
M_MN249 N$296 N$297 0 0 n l=2e-06 w=6e-06
M_MN547 N$11786 RST 0 0 n l=2e-06 w=5e-06
M_MN140 N$158 N$389 0 0 n l=2e-06 w=3e-06
M_MN401 N$11804 N$1674 N$11805 0 n l=2e-06 w=3e-06
M_MN451 N$1615 N$1620 0 0 n l=2e-06 w=3e-06
M_MN450 N$9715 N$1633 N$1616 0 n l=2e-06 w=3e-06
M_MN449 N$1616 N$1599 0 0 n l=2e-06 w=3e-06
M_MN448 N$13447 N$9715 0 0 n l=2e-06 w=3e-06
M_MN242 N$283 CK 0 0 n l=2e-06 w=5e-06
M_MN68 N$290 N$288 0 0 n l=2e-06 w=6e-06
M_MN272 N$315 N$312 0 0 n l=2e-06 w=6e-06
M_MN303 N$338 N$339 0 0 n l=2e-06 w=6e-06
M_MN279 N$319 N$320 N$254 0 n l=2e-06 w=6e-06
M_MN278 N$313 CK 0 0 n l=2e-06 w=5e-06
M_MN283 N$323 CK N$321 0 n l=2e-06 w=6e-06
M_MN250 N$297 N$295 0 0 n l=2e-06 w=6e-06
M_MN220 N$254 N$265 N$200 0 n l=2e-06 w=5e-06
M_MN219 N$254 N$14095 N$183 0 n l=2e-06 w=5e-06
M_MN280 N$321 CK N$319 0 n l=2e-06 w=6e-06
M_MN286 N$325 N$323 0 0 n l=2e-06 w=6e-06
M_MN226 N$262 N$265 N$1179 0 n l=2e-06 w=5e-06
M_MN225 N$262 N$14095 N$217 0 n l=2e-06 w=5e-06
M_MN67 N$361 N$290 0 0 n l=2e-06 w=6e-06
M_MN526 N$1558 N$1551 N$1547 0 n l=2e-06 w=6e-06
M_MN213 N$246 N$14095 N$148 0 n l=2e-06 w=5e-06
M_MN256 N$302 CK N$300 0 n l=2e-06 w=6e-06
M_MN255 N$300 N$301 0 0 n l=2e-06 w=6e-06
M_MN139 N$154 N$138 N$157 0 n l=2e-06 w=3e-06
M_MN168 N$192 N$392 0 0 n l=2e-06 w=3e-06
M_MN167 N$188 N$173 N$191 0 n l=2e-06 w=3e-06
M_MN166 N$191 N$14079 0 0 n l=2e-06 w=3e-06
M_MN165 N$190 N$188 0 0 n l=2e-06 w=3e-06
M_MN318 N$14084 N$11347 0 0 n l=2e-06 w=5e-06
M_MN317 N$348 N$11347 0 0 n l=2e-06 w=5e-06
M_MN316 OUT8 N$348 N$361 0 n l=2e-06 w=5e-06
M_MN331 N$14090 N$11347 0 0 n l=2e-06 w=5e-06
M_MN769 N$11802 C N$11804 0 n l=2e-06 w=3e-06
M_MN400 N$11803 C 0 0 n l=2e-06 w=3e-06
M_MN399 N$11803 N$11794 0 0 n l=2e-06 w=3e-06
M_MN398 N$11803 N$1674 0 0 n l=2e-06 w=3e-06
M_MN459 N$1611 N$9715 N$1610 0 n l=2e-06 w=3e-06
M_MN458 N$1608 N$1620 0 0 n l=2e-06 w=3e-06
M_MN464 N$1620 0 0 0 n l=2e-06 w=3e-06
M_MN351 N$396 N$14095 N$14091 0 n l=2e-06 w=5e-06
M_MN731 N$11099 N$11321 N$11324 0 n l=2e-06 w=6e-06
M_MN721 N$11318 CK N$11316 0 n l=2e-06 w=6e-06
M_MN720 N$11316 N$11317 0 0 n l=2e-06 w=6e-06
M_MN719 N$11317 N$11314 0 0 n l=2e-06 w=6e-06
M_MN718 N$11316 CK N$11314 0 n l=2e-06 w=6e-06
M_MN752 N$11336 CK N$11334 0 n l=2e-06 w=6e-06
M_MN753 N$382 N$11333 N$11336 0 n l=2e-06 w=6e-06
M_MN352 N$396 N$11347 N$345 0 n l=2e-06 w=5e-06
M_MN535 N$1554 N$1544 N$1540 0 n l=2e-06 w=6e-06
M_MN534 N$1540 CK N$1542 0 n l=2e-06 w=6e-06
M_MN887 N$14029 N$14037 P3 0 n l=2e-06 w=5e-06
M_MN895 N$14024 SK1 0 0 n l=2e-06 w=5e-06
M_MN525 N$1547 CK N$1549 0 n l=2e-06 w=6e-06
M_MN524 N$1549 N$1548 0 0 n l=2e-06 w=6e-06
M_MN530 N$1545 N$1544 N$13447 0 n l=2e-06 w=6e-06
M_MN529 N$1551 CK 0 0 n l=2e-06 w=6e-06
M_MN528 N$1546 N$1547 0 0 n l=2e-06 w=6e-06
M_MN527 N$1558 N$1546 0 0 n l=2e-06 w=6e-06
M_MN533 N$1542 N$1541 0 0 n l=2e-06 w=6e-06
M_MN548 N$11786 N$11813 N$12632 0 n l=2e-06 w=5e-06
M_MN482 N$1585 CK N$1589 0 n l=2e-06 w=6e-06
M_MN481 N$1589 N$1588 N$1593 0 n l=2e-06 w=6e-06
M_MN480 N$1593 N$13243 N$1674 0 n l=2e-06 w=5e-06
M_MN877 N$14039 N$14040 0 0 n l=2e-06 w=5e-06
M_MN888 N$14029 N$14040 0 0 n l=2e-06 w=5e-06
M_MN876 N$14039 N$14037 0 0 n l=2e-06 w=5e-06
M_MN906 N$14018 N$14024 N$14028 0 n l=2e-06 w=5e-06
M_MN911 N$14016 SK2 N$14022 0 n l=2e-06 w=5e-06
M_MN463 N$1653 B2 0 0 n l=2e-06 w=3e-06
M_MN462 N$1673 B1 0 0 n l=2e-06 w=3e-06
M_MN460 N$1611 N$1633 N$1609 0 n l=2e-06 w=3e-06
M_MN466 N$13650 N$11810 0 0 n l=2e-06 w=6e-06
M_MN465 N$1636 B3 0 0 n l=2e-06 w=3e-06
M_MN540 N$1674 RST A5 0 n l=2e-06 w=5e-06
M_MN884 N$14031 N$14040 0 0 n l=2e-06 w=5e-06
M_MN889 N$14028 N$14037 P2 0 n l=2e-06 w=5e-06
M_MN376 N$11790 CK N$11783 0 n l=2e-06 w=6e-06
M_MN375 N$11783 N$11782 0 0 n l=2e-06 w=6e-06
M_MN381 N$11781 N$11780 N$11817 0 n l=2e-06 w=6e-06
M_MN380 N$11789 CK 0 0 n l=2e-06 w=5e-06
M_MN894 N$14025 SK1 N$14035 0 n l=2e-06 w=5e-06
M_MN893 N$14025 N$14024 N$14039 0 n l=2e-06 w=5e-06
M_MN898 N$14022 N$14024 N$14033 0 n l=2e-06 w=5e-06
M_MN897 N$14023 SK1 N$14033 0 n l=2e-06 w=5e-06
M_MN896 N$14023 N$14024 N$14035 0 n l=2e-06 w=5e-06
M_MN901 N$14021 SK1 N$14030 0 n l=2e-06 w=5e-06
M_MN934 N$14003 N$14006 N$14012 0 n l=2e-06 w=5e-06
M_MN940 N$14000 N$14006 N$14009 0 n l=2e-06 w=5e-06
M_MN939 N$14001 SK3 0 0 n l=2e-06 w=5e-06
M_MN741 N$11088 N$11331 0 0 n l=2e-06 w=6e-06
M_MN743 N$11327 CK 0 0 n l=2e-06 w=5e-06
M_MN361 N$388 N$409 N$374 0 n l=2e-06 w=5e-06
M_MN2 N$6 N$3 0 0 n l=2e-06 w=6e-06
M_MN910 N$14016 N$14015 N$14025 0 n l=2e-06 w=5e-06
M_MN909 N$14017 SK1 0 0 n l=2e-06 w=5e-06
M_MN914 N$14014 SK2 N$14021 0 n l=2e-06 w=5e-06
M_MN913 N$14014 N$14015 N$14023 0 n l=2e-06 w=5e-06
M_MN912 N$14015 SK2 0 0 n l=2e-06 w=5e-06
M_MN917 N$14012 N$14015 N$14021 0 n l=2e-06 w=5e-06
M_MN881 N$14033 N$14037 0 0 n l=2e-06 w=5e-06
M_MN886 N$14030 N$14040 0 0 n l=2e-06 w=5e-06
M_MN885 N$14030 N$14037 P4 0 n l=2e-06 w=5e-06
M_MN16 N$24 N$22 0 0 n l=2e-06 w=6e-06
M_MN21 N$27 N$14 N$29 0 n l=2e-06 w=6e-06
M_MN229 N$266 N$265 N$1180 0 n l=2e-06 w=5e-06
M_MN324 N$14087 N$11347 0 0 n l=2e-06 w=5e-06
M_MN356 N$386 N$14096 P1 0 n l=2e-06 w=5e-06
M_MN6 N$12 N$10 0 0 n l=2e-06 w=6e-06
M_MN5 N$8 N$3 N$12 0 n l=2e-06 w=6e-06
M_MN4 N$11 add_one 0 0 n l=2e-06 w=6e-06
M_MN3 N$8 N$9 N$11 0 n l=2e-06 w=6e-06
M_MN379 N$11787 N$11790 0 0 n l=2e-06 w=6e-06
M_MN384 N$11779 N$11778 0 0 n l=2e-06 w=6e-06
M_MN383 N$11778 N$11781 0 0 n l=2e-06 w=6e-06
M_MN892 N$14027 N$14040 0 0 n l=2e-06 w=5e-06
M_MN891 N$14027 N$14037 P1 0 n l=2e-06 w=5e-06
M_MN932 N$14004 N$14006 N$14013 0 n l=2e-06 w=5e-06
M_MN931 N$14005 SK3 N$14011 0 n l=2e-06 w=5e-06
M_MN937 N$14002 SK3 N$14008 0 n l=2e-06 w=5e-06
M_MN936 N$14002 N$14006 N$14011 0 n l=2e-06 w=5e-06
M_MN935 N$14003 SK3 N$14009 0 n l=2e-06 w=5e-06
M_MN9 N$13 N$8 0 0 n l=2e-06 w=6e-06
M_MN8 N$10 add_one 0 0 n l=2e-06 w=6e-06
M_MN505 N$12429 N$12633 0 0 n l=2e-06 w=6e-06
M_MN404 N$1177 0 0 0 n l=2e-06 w=5e-06
M_MN591 SK3 N$1491 0 0 n l=2e-06 w=6e-06
M_MN1 N$2 add_one N$6 0 n l=2e-06 w=6e-06
M_MN241 N$279 N$385 0 0 n l=2e-06 w=6e-06
M_MN742 N$11331 N$11330 0 0 n l=2e-06 w=6e-06
M_MN405 N$1180 N$1177 0 0 n l=2e-06 w=5e-06
M_MN323 N$14086 N$348 N$310 0 n l=2e-06 w=5e-06
M_MN325 N$14087 N$348 N$317 0 n l=2e-06 w=5e-06
M_MN18 N$22 N$17 0 0 n l=2e-06 w=6e-06
M_MN17 N$21 N$16 0 0 n l=2e-06 w=6e-06
M_MN252 N$298 N$299 N$242 0 n l=2e-06 w=6e-06
M_MN150 N$166 N$162 0 0 n l=2e-06 w=3e-06
M_MN149 N$162 N$138 N$164 0 n l=2e-06 w=3e-06
M_MN148 N$162 N$154 N$163 0 n l=2e-06 w=3e-06
M_MN117 N$127 N$102 0 0 n l=2e-06 w=3e-06
M_MN116 N$127 N$387 0 0 n l=2e-06 w=3e-06
M_MN368 N$394 N$14096 0 0 n l=2e-06 w=5e-06
M_MN367 N$392 N$409 N$412 0 n l=2e-06 w=5e-06
M_MN366 N$392 N$14096 0 0 n l=2e-06 w=5e-06
M_MN452 N$1616 N$1620 0 0 n l=2e-06 w=3e-06
M_MN447 N$12835 N$1627 0 0 n l=2e-06 w=3e-06
M_MN446 N$1627 N$1650 N$1625 0 n l=2e-06 w=3e-06
M_MN61 N$282 N$283 N$271 0 n l=2e-06 w=6e-06
M_MN228 N$266 N$14095 N$1179 0 n l=2e-06 w=5e-06
M_MN345 N$376 N$14095 N$14088 0 n l=2e-06 w=5e-06
M_MN371 N$395 N$409 N$396 0 n l=2e-06 w=5e-06
M_MN305 N$334 CK 0 0 n l=2e-06 w=5e-06
M_MN304 N$339 N$337 0 0 n l=2e-06 w=6e-06
M_MN314 N$341 CK 0 0 n l=2e-06 w=5e-06
M_MN98 N$104 N$386 0 0 n l=2e-06 w=3e-06
M_MN127 N$139 N$388 0 0 n l=2e-06 w=3e-06
M_MN267 N$310 N$311 0 0 n l=2e-06 w=6e-06
M_MN748 N$11332 N$11333 N$11083 0 n l=2e-06 w=6e-06
M_MN403 N$1177 N$1179 0 0 n l=2e-06 w=5e-06
M_MN268 N$311 N$309 0 0 n l=2e-06 w=6e-06
M_MN369 N$394 N$409 N$397 0 n l=2e-06 w=5e-06
M_MN326 N$14091 N$11347 0 0 n l=2e-06 w=5e-06
M_MN348 N$412 N$11347 N$331 0 n l=2e-06 w=5e-06
M_MN311 N$345 N$341 N$344 0 n l=2e-06 w=6e-06
M_MN178 N$200 N$196 0 0 n l=2e-06 w=3e-06
M_MN132 N$146 0 N$147 0 n l=2e-06 w=3e-06
M_MN131 N$145 N$120 0 0 n l=2e-06 w=3e-06
M_MN129 N$145 0 0 0 n l=2e-06 w=3e-06
M_MN773 N$1599 N$11813 N$12429 0 n l=2e-06 w=5e-06
M_MN294 N$331 N$332 0 0 n l=2e-06 w=6e-06
M_MN772 N$1599 RST 0 0 n l=2e-06 w=5e-06
M_MN771 N$11794 B0 0 0 n l=2e-06 w=3e-06
M_MN485 N$1583 CK N$1585 0 n l=2e-06 w=6e-06
M_MN484 N$1585 N$1584 0 0 n l=2e-06 w=6e-06
M_MN354 N$385 N$409 N$398 0 n l=2e-06 w=5e-06
M_MN353 N$385 N$14096 0 0 n l=2e-06 w=5e-06
M_MN343 N$411 N$14095 N$14087 0 n l=2e-06 w=5e-06
M_MN313 N$346 N$344 0 0 n l=2e-06 w=6e-06
M_MN192 N$217 N$213 0 0 n l=2e-06 w=3e-06
M_MN147 N$165 N$389 0 0 n l=2e-06 w=3e-06
M_MN146 N$164 0 N$165 0 n l=2e-06 w=3e-06
M_MN115 N$127 0 0 0 n l=2e-06 w=3e-06
M_MN144 N$163 N$389 0 0 n l=2e-06 w=3e-06
M_MN143 N$163 0 0 0 n l=2e-06 w=3e-06
M_MN199 N$231 N$14081 0 0 n l=2e-06 w=3e-06
M_MN126 N$140 N$388 0 0 n l=2e-06 w=3e-06
M_MN125 N$136 N$120 N$139 0 n l=2e-06 w=3e-06
M_MN124 N$139 0 0 0 n l=2e-06 w=3e-06
M_MN153 N$171 N$156 N$174 0 n l=2e-06 w=3e-06
M_MN152 N$174 N$14078 0 0 n l=2e-06 w=3e-06
M_MN151 N$173 N$171 0 0 n l=2e-06 w=3e-06
M_MN284 N$324 N$320 N$323 0 n l=2e-06 w=6e-06
M_MN62 N$286 CK N$282 0 n l=2e-06 w=6e-06
M_MN66 N$361 N$283 N$288 0 n l=2e-06 w=6e-06
M_MN285 N$324 N$325 0 0 n l=2e-06 w=6e-06
M_MN689 N$14098 CK 0 0 n l=2e-06 w=5e-06
M_MN643 N$1441 N$1462 N$1439 0 n l=2e-06 w=3e-06
M_MN642 N$1441 N$1448 N$1440 0 n l=2e-06 w=3e-06
M_MN641 N$1438 N$1450 0 0 n l=2e-06 w=3e-06
M_MN647 N$1433 N$1447 N$1431 0 n l=2e-06 w=3e-06
M_MN646 N$1431 B3 0 0 n l=2e-06 w=3e-06
M_MN675 N$1410 N$1557 N$1452 0 n l=2e-06 w=5e-06
M_MN681 N$1406 N$14098 N$14097 0 n l=2e-06 w=6e-06
M_MN254 N$301 N$298 0 0 n l=2e-06 w=6e-06
M_MN302 N$338 N$334 N$337 0 n l=2e-06 w=6e-06
M_MN301 N$337 CK N$335 0 n l=2e-06 w=6e-06
M_MN300 N$335 N$336 0 0 n l=2e-06 w=6e-06
M_MN251 N$292 CK 0 0 n l=2e-06 w=5e-06
M_MN232 N$271 N$265 N$112 0 n l=2e-06 w=5e-06
M_MN847 OUT5 N$13959 0 0 n l=2e-06 w=3e-06
M_MN875 OUT7 N$13991 0 0 n l=2e-06 w=3e-06
M_MN874 N$13991 N$13969 N$13993 0 n l=2e-06 w=3e-06
M_MN710 N$1385 N$1388 0 0 n l=2e-06 w=6e-06
M_MN177 N$196 N$173 N$198 0 n l=2e-06 w=3e-06
M_MN716 N$1387 CK 0 0 n l=2e-06 w=5e-06
M_MN686 N$14046 N$14098 N$1402 0 n l=2e-06 w=6e-06
M_MN685 N$1402 CK N$1404 0 n l=2e-06 w=6e-06
M_MN691 N$1398 CK N$1400 0 n l=2e-06 w=6e-06
M_MN690 N$1400 N$1399 N$1410 0 n l=2e-06 w=6e-06
M_MN163 N$179 N$156 N$181 0 n l=2e-06 w=3e-06
M_MN162 N$179 N$171 N$180 0 n l=2e-06 w=3e-06
M_MN295 N$332 N$330 0 0 n l=2e-06 w=6e-06
M_MN680 N$1408 N$1413 0 0 n l=2e-06 w=5e-06
M_MN679 N$1408 N$1557 N$1422 0 n l=2e-06 w=5e-06
M_MN880 N$14035 N$14040 0 0 n l=2e-06 w=5e-06
M_MN879 N$14035 N$14037 0 0 n l=2e-06 w=5e-06
M_MN878 N$14037 N$14040 0 0 n l=2e-06 w=5e-06
M_MN883 N$14031 N$14037 0 0 n l=2e-06 w=5e-06
M_MN882 N$14033 N$14040 0 0 n l=2e-06 w=5e-06
M_MN873 N$13991 N$13983 N$13992 0 n l=2e-06 w=3e-06
M_MN751 N$11334 N$11335 0 0 n l=2e-06 w=6e-06
M_MN750 N$11335 N$11332 0 0 n l=2e-06 w=6e-06
M_MN736 N$11328 CK N$11326 0 n l=2e-06 w=6e-06
M_MN735 N$11326 N$11327 N$11344 0 n l=2e-06 w=6e-06
M_MN734 N$11321 CK 0 0 n l=2e-06 w=5e-06
M_MN733 N$11325 N$11324 0 0 n l=2e-06 w=6e-06
M_MN732 N$11099 N$11325 0 0 n l=2e-06 w=6e-06
M_MN359 N$387 N$409 N$410 0 n l=2e-06 w=5e-06
M_MN360 N$388 N$14096 P3 0 n l=2e-06 w=5e-06
M_MN164 N$183 N$179 0 0 n l=2e-06 w=3e-06
M_MP106 N$108 N$84 N$107 VDD p l=2e-06 w=3e-06
M_MP105 N$107 N$386 N$106 VDD p l=2e-06 w=3e-06
M_MP104 N$106 0 N$105 VDD p l=2e-06 w=3e-06
M_MP103 N$105 N$386 VDD VDD p l=2e-06 w=3e-06
M_MP102 N$105 0 VDD VDD p l=2e-06 w=3e-06
M_MP146 N$160 0 N$159 VDD p l=2e-06 w=3e-06
M_MP145 N$159 N$389 VDD VDD p l=2e-06 w=3e-06
M_MP144 N$159 0 VDD VDD p l=2e-06 w=3e-06
M_MP143 N$159 N$138 VDD VDD p l=2e-06 w=3e-06
M_MP187 N$210 N$394 VDD VDD p l=2e-06 w=3e-06
M_MP253 N$298 N$299 N$300 VDD p l=2e-06 w=6e-06
M_MP294 N$331 N$332 VDD VDD p l=2e-06 w=6e-06
M_MP293 N$330 CK N$331 VDD p l=2e-06 w=6e-06
M_MP292 N$328 N$327 N$330 VDD p l=2e-06 w=6e-06
M_MP345 N$14088 N$11347 N$376 VDD p l=2e-06 w=5e-06
M_MP16 N$20 N$17 N$19 VDD p l=2e-06 w=6e-06
M_MP356 P1 N$409 N$386 VDD p l=2e-06 w=5e-06
M_MP391 0 N$13447 N$11570 VDD p l=2e-06 w=5e-06
M_MP390 N$1674 N$13243 N$11570 VDD p l=2e-06 w=5e-06
M_MP55 N$25 N$419 N$61 VDD p l=2e-06 w=6e-06
M_MP54 0 N$420 N$60 VDD p l=2e-06 w=6e-06
M_MP59 N$46 N$419 N$63 VDD p l=2e-06 w=6e-06
M_MP58 0 N$420 N$62 VDD p l=2e-06 w=6e-06
M_MP71 N$66 N$65 VDD VDD p l=2e-06 w=5e-06
M_MP77 N$72 N$71 VDD VDD p l=2e-06 w=5e-06
M_MP76 N$71 N$61 N$70 VDD p l=2e-06 w=5e-06
M_MP75 N$70 N$60 VDD VDD p l=2e-06 w=5e-06
M_MP80 N$75 N$74 VDD VDD p l=2e-06 w=5e-06
M_MP79 N$74 N$63 N$73 VDD p l=2e-06 w=5e-06
M_MP78 N$73 N$62 VDD VDD p l=2e-06 w=5e-06
M_MP951 N$14074 N$11345 VDD VDD p l=2e-06 w=5e-06
M_MP950 N$66 N$11345 N$14078 VDD p l=2e-06 w=5e-06
M_MP949 0 N$14074 N$14078 VDD p l=2e-06 w=5e-06
M_MP957 N$75 N$11345 N$14081 VDD p l=2e-06 w=5e-06
M_MP44 N$16 N$14093 VDD VDD p l=2e-06 w=6e-06
M_MP43 N$3 N$14046 VDD VDD p l=2e-06 w=6e-06
M_MP42 N$38 N$14092 VDD VDD p l=2e-06 w=6e-06
M_MP47 N$13 N$419 N$56 VDD p l=2e-06 w=6e-06
M_MP46 0 N$420 N$53 VDD p l=2e-06 w=6e-06
M_MP956 0 N$14074 N$14081 VDD p l=2e-06 w=5e-06
M_MP955 N$72 N$11345 N$14080 VDD p l=2e-06 w=5e-06
M_MP954 0 N$14074 N$14080 VDD p l=2e-06 w=5e-06
M_MP953 N$415 N$11345 N$14079 VDD p l=2e-06 w=5e-06
M_MP952 0 N$14074 N$14079 VDD p l=2e-06 w=5e-06
M_MP53 N$14093 N$417 N$60 VDD p l=2e-06 w=6e-06
M_MP52 0 N$421 N$59 VDD p l=2e-06 w=6e-06
M_MP51 N$36 N$419 N$59 VDD p l=2e-06 w=6e-06
M_MP50 0 N$420 N$58 VDD p l=2e-06 w=6e-06
M_MP57 N$14092 N$417 N$62 VDD p l=2e-06 w=6e-06
M_MP56 0 N$421 N$61 VDD p l=2e-06 w=6e-06
M_MP28 N$33 N$14 VDD VDD p l=2e-06 w=6e-06
M_MP27 N$32 N$28 VDD VDD p l=2e-06 w=6e-06
M_MP32 N$37 N$26 VDD VDD p l=2e-06 w=6e-06
M_MP31 N$37 N$38 VDD VDD p l=2e-06 w=6e-06
M_MP70 N$65 N$56 N$64 VDD p l=2e-06 w=5e-06
M_MP69 N$64 N$53 VDD VDD p l=2e-06 w=5e-06
M_MP60 0 N$421 N$63 VDD p l=2e-06 w=6e-06
M_MP74 N$415 N$68 VDD VDD p l=2e-06 w=5e-06
M_MP73 N$68 N$59 N$67 VDD p l=2e-06 w=5e-06
M_MP72 N$67 N$58 VDD VDD p l=2e-06 w=5e-06
M_MP37 N$42 N$38 VDD VDD p l=2e-06 w=6e-06
M_MP41 N$28 N$14045 VDD VDD p l=2e-06 w=6e-06
M_MP40 H_A_Cout N$37 VDD VDD p l=2e-06 w=6e-06
M_MP39 N$46 N$41 VDD VDD p l=2e-06 w=6e-06
M_MP365 N$376 N$14096 N$390 VDD p l=2e-06 w=5e-06
M_MP364 0 N$409 N$390 VDD p l=2e-06 w=5e-06
M_MP363 N$411 N$14096 N$389 VDD p l=2e-06 w=5e-06
M_MP362 P4 N$409 N$389 VDD p l=2e-06 w=5e-06
M_MP97 N$99 N$386 N$96 VDD p l=2e-06 w=3e-06
M_MP5 N$7 N$10 VDD VDD p l=2e-06 w=6e-06
M_MP4 N$8 N$9 N$7 VDD p l=2e-06 w=6e-06
M_MP3 N$7 N$3 VDD VDD p l=2e-06 w=6e-06
M_MP45 N$14046 N$417 N$53 VDD p l=2e-06 w=6e-06
M_MP49 N$14045 N$417 N$58 VDD p l=2e-06 w=6e-06
M_MP48 0 N$421 N$56 VDD p l=2e-06 w=6e-06
M_MP22 N$27 N$14 VDD VDD p l=2e-06 w=6e-06
M_MP21 N$27 N$28 VDD VDD p l=2e-06 w=6e-06
M_MP20 N$26 N$15 VDD VDD p l=2e-06 w=6e-06
M_MP26 N$31 N$14 N$30 VDD p l=2e-06 w=6e-06
M_MP25 N$30 N$33 VDD VDD p l=2e-06 w=6e-06
M_MP24 N$31 N$32 N$30 VDD p l=2e-06 w=6e-06
M_MP23 N$30 N$28 VDD VDD p l=2e-06 w=6e-06
M_MP335 N$361 N$14095 N$398 VDD p l=2e-06 w=5e-06
M_MP371 N$396 N$14096 N$395 VDD p l=2e-06 w=5e-06
M_MP7 N$9 N$3 VDD VDD p l=2e-06 w=6e-06
M_MP30 N$17 N$27 VDD VDD p l=2e-06 w=6e-06
M_MP29 N$36 N$31 VDD VDD p l=2e-06 w=6e-06
M_MP36 N$41 N$26 N$40 VDD p l=2e-06 w=6e-06
M_MP35 N$40 N$43 VDD VDD p l=2e-06 w=6e-06
M_MP34 N$41 N$42 N$40 VDD p l=2e-06 w=6e-06
M_MP33 N$40 N$38 VDD VDD p l=2e-06 w=6e-06
M_MP38 N$43 N$26 VDD VDD p l=2e-06 w=6e-06
M_MP324 0 N$348 N$14087 VDD p l=2e-06 w=5e-06
M_MP325 N$317 N$11347 N$14087 VDD p l=2e-06 w=5e-06
M_MP739 N$11328 N$11327 N$11330 VDD p l=2e-06 w=6e-06
M_MP767 N$11347 N$11345 VDD VDD p l=2e-06 w=5e-06
M_MP727 N$11320 N$11321 N$11322 VDD p l=2e-06 w=6e-06
M_MP726 N$14096 CK N$11320 VDD p l=2e-06 w=6e-06
M_MP725 N$11315 CK VDD VDD p l=2e-06 w=5e-06
M_MP82 N$77 N$385 VDD VDD p l=2e-06 w=3e-06
M_MP81 N$77 0 VDD VDD p l=2e-06 w=3e-06
M_MP740 N$11330 CK N$11088 VDD p l=2e-06 w=6e-06
M_MP271 N$312 N$313 N$314 VDD p l=2e-06 w=6e-06
M_MP270 N$250 CK N$312 VDD p l=2e-06 w=6e-06
M_MP737 N$11329 N$11326 VDD VDD p l=2e-06 w=6e-06
M_MP736 N$11326 N$11327 N$11328 VDD p l=2e-06 w=6e-06
M_MP741 N$11088 N$11331 VDD VDD p l=2e-06 w=6e-06
M_MP350 N$338 N$14095 N$397 VDD p l=2e-06 w=5e-06
M_MP338 N$296 N$14095 N$372 VDD p l=2e-06 w=5e-06
M_MP337 N$14084 N$11347 N$372 VDD p l=2e-06 w=5e-06
M_MP336 N$14095 N$11347 VDD VDD p l=2e-06 w=5e-06
M_MP11 N$15 N$16 VDD VDD p l=2e-06 w=6e-06
M_MP383 N$11778 N$11781 VDD VDD p l=2e-06 w=6e-06
M_MP382 N$11781 N$11780 N$11779 VDD p l=2e-06 w=6e-06
M_MP388 N$11775 N$11777 VDD VDD p l=2e-06 w=6e-06
M_MP387 N$12632 N$11775 VDD VDD p l=2e-06 w=6e-06
M_MP386 N$11777 CK N$12632 VDD p l=2e-06 w=6e-06
M_MP385 N$11779 N$11780 N$11777 VDD p l=2e-06 w=6e-06
M_MP322 0 N$348 N$14086 VDD p l=2e-06 w=5e-06
M_MP321 N$384 N$11347 N$14085 VDD p l=2e-06 w=5e-06
M_MP158 N$176 N$14078 VDD VDD p l=2e-06 w=3e-06
M_MP157 N$176 N$156 VDD VDD p l=2e-06 w=3e-06
M_MP186 N$210 N$14080 VDD VDD p l=2e-06 w=3e-06
M_MP361 N$374 N$14096 N$388 VDD p l=2e-06 w=5e-06
M_MP191 N$213 N$205 N$210 VDD p l=2e-06 w=3e-06
M_MP190 N$213 N$190 N$212 VDD p l=2e-06 w=3e-06
M_MP189 N$212 N$394 N$211 VDD p l=2e-06 w=3e-06
M_MP188 N$211 N$14080 N$210 VDD p l=2e-06 w=3e-06
M_MP213 N$148 N$265 N$246 VDD p l=2e-06 w=5e-06
M_MP729 N$11322 N$11323 VDD VDD p l=2e-06 w=6e-06
M_MP728 N$11323 N$11320 VDD VDD p l=2e-06 w=6e-06
M_MP328 N$324 N$11347 N$14088 VDD p l=2e-06 w=5e-06
M_MP327 0 N$348 N$14088 VDD p l=2e-06 w=5e-06
M_MP326 0 N$348 N$14091 VDD p l=2e-06 w=5e-06
M_MP332 N$338 N$11347 N$14090 VDD p l=2e-06 w=5e-06
M_MP183 N$205 N$14080 N$204 VDD p l=2e-06 w=3e-06
M_MP182 N$205 N$190 N$202 VDD p l=2e-06 w=3e-06
M_MP330 N$331 N$11347 N$14089 VDD p l=2e-06 w=5e-06
M_MP297 N$262 CK N$333 VDD p l=2e-06 w=6e-06
M_MP723 N$14096 N$11319 VDD VDD p l=2e-06 w=6e-06
M_MP722 N$11318 CK N$14096 VDD p l=2e-06 w=6e-06
M_MP747 N$11108 N$11344 N$11104 VDD p l=2e-06 w=5e-06
M_MP746 N$11104 N$11099 N$11100 VDD p l=2e-06 w=5e-06
M_MP745 N$11100 N$14096 N$11096 VDD p l=2e-06 w=5e-06
M_MP744 N$11096 N$382 VDD VDD p l=2e-06 w=5e-06
M_MP749 N$11332 N$11333 N$11334 VDD p l=2e-06 w=6e-06
M_MP748 N$11083 CK N$11332 VDD p l=2e-06 w=6e-06
M_MP378 N$14107 N$11787 VDD VDD p l=2e-06 w=6e-06
M_MP663 N$1488 N$1416 N$1521 VDD p l=2e-06 w=5e-06
M_MP662 N$1450 N$1485 VDD VDD p l=2e-06 w=3e-06
M_MP693 N$1398 N$1397 VDD VDD p l=2e-06 w=6e-06
M_MP702 N$1392 N$1391 VDD VDD p l=2e-06 w=6e-06
M_MP701 N$1391 N$1394 VDD VDD p l=2e-06 w=6e-06
M_MP707 N$1393 CK VDD VDD p l=2e-06 w=5e-06
M_MP706 N$1389 N$1390 VDD VDD p l=2e-06 w=6e-06
M_MP705 N$14093 N$1389 VDD VDD p l=2e-06 w=6e-06
M_MP704 N$1390 CK N$14093 VDD p l=2e-06 w=6e-06
M_MP342 N$310 N$14095 N$374 VDD p l=2e-06 w=5e-06
M_MP341 N$14086 N$11347 N$374 VDD p l=2e-06 w=5e-06
M_MP141 N$154 0 N$153 VDD p l=2e-06 w=3e-06
M_MP140 N$154 N$138 N$150 VDD p l=2e-06 w=3e-06
M_MP139 N$153 N$389 N$150 VDD p l=2e-06 w=3e-06
M_MP696 N$14045 N$1395 VDD VDD p l=2e-06 w=6e-06
M_MP695 N$1396 CK N$14045 VDD p l=2e-06 w=6e-06
M_MP694 N$1398 N$1399 N$1396 VDD p l=2e-06 w=6e-06
M_MP700 N$1394 N$1393 N$1392 VDD p l=2e-06 w=6e-06
M_MP659 N$1481 N$1488 VDD VDD p l=2e-06 w=3e-06
M_MP660 N$1465 N$1486 VDD VDD p l=2e-06 w=3e-06
M_MP708 N$1408 CK N$1388 VDD p l=2e-06 w=6e-06
M_MP730 N$11322 N$11321 N$11324 VDD p l=2e-06 w=6e-06
M_MP85 N$81 0 N$80 VDD p l=2e-06 w=3e-06
M_MP84 N$81 0 N$77 VDD p l=2e-06 w=3e-06
M_MP673 0 N$1557 N$14097 VDD p l=2e-06 w=5e-06
M_MP15 N$19 N$22 VDD VDD p l=2e-06 w=6e-06
M_MP14 N$20 N$21 N$19 VDD p l=2e-06 w=6e-06
M_MP13 N$19 N$16 VDD VDD p l=2e-06 w=6e-06
M_MP891 P1 N$14040 N$14027 VDD p l=2e-06 w=5e-06
M_MP343 N$14087 N$11347 N$411 VDD p l=2e-06 w=5e-06
M_MP738 N$11328 N$11329 VDD VDD p l=2e-06 w=6e-06
M_MP313 N$346 N$344 VDD VDD p l=2e-06 w=6e-06
M_MP312 N$345 N$346 VDD VDD p l=2e-06 w=6e-06
M_MP127 N$136 0 N$135 VDD p l=2e-06 w=3e-06
M_MP126 N$136 N$120 N$132 VDD p l=2e-06 w=3e-06
M_MP125 N$135 N$388 N$132 VDD p l=2e-06 w=3e-06
M_MP710 N$1385 N$1388 VDD VDD p l=2e-06 w=6e-06
M_MP709 N$1388 N$1387 N$1386 VDD p l=2e-06 w=6e-06
M_MP296 N$327 CK VDD VDD p l=2e-06 w=5e-06
M_MP542 N$11813 RST VDD VDD p l=2e-06 w=5e-06
M_MP574 N$1507 N$1509 VDD VDD p l=2e-06 w=6e-06
M_MP551 N$1530 N$14108 VDD VDD p l=2e-06 w=5e-06
M_MP550 0 N$14108 N$1529 VDD p l=2e-06 w=5e-06
M_MP549 N$14107 N$1530 N$1529 VDD p l=2e-06 w=5e-06
M_MP666 N$1486 N$1416 N$1512 VDD p l=2e-06 w=5e-06
M_MP691 N$1400 N$1399 N$1398 VDD p l=2e-06 w=6e-06
M_MP697 N$1395 N$1396 VDD VDD p l=2e-06 w=6e-06
M_MP424 N$1651 N$11561 N$1652 VDD p l=2e-06 w=3e-06
M_MP423 N$1651 N$1668 N$1655 VDD p l=2e-06 w=3e-06
M_MP428 N$1647 N$1653 VDD VDD p l=2e-06 w=3e-06
M_MP427 N$1647 N$11561 VDD VDD p l=2e-06 w=3e-06
M_MP538 N$1544 CK VDD VDD p l=2e-06 w=5e-06
M_MP765 N$11339 CK VDD VDD p l=2e-06 w=5e-06
M_MP703 N$1392 N$1393 N$1390 VDD p l=2e-06 w=6e-06
M_MP670 N$1484 N$1416 N$1496 VDD p l=2e-06 w=5e-06
M_MP675 N$1452 N$1413 N$1410 VDD p l=2e-06 w=5e-06
M_MP674 N$1413 N$1557 VDD VDD p l=2e-06 w=5e-06
M_MP759 N$11341 N$11338 VDD VDD p l=2e-06 w=6e-06
M_MP758 N$11338 N$11339 N$11340 VDD p l=2e-06 w=6e-06
M_MP757 N$11099 CK N$11338 VDD p l=2e-06 w=6e-06
M_MP756 N$11333 CK VDD VDD p l=2e-06 w=5e-06
M_MP755 N$11337 N$11336 VDD VDD p l=2e-06 w=6e-06
M_MP770 N$11810 N$11802 VDD VDD p l=2e-06 w=3e-06
M_MP520 N$13857 N$1558 VDD VDD p l=2e-06 w=5e-06
M_MP519 N$13857 N$1554 VDD VDD p l=2e-06 w=5e-06
M_MP724 N$11319 N$11318 VDD VDD p l=2e-06 w=6e-06
M_MP124 N$132 N$388 VDD VDD p l=2e-06 w=3e-06
M_MP315 0 N$348 OUT8 VDD p l=2e-06 w=5e-06
M_MP295 N$332 N$330 VDD VDD p l=2e-06 w=6e-06
M_MP349 N$14090 N$11347 N$397 VDD p l=2e-06 w=5e-06
M_MP348 N$331 N$14095 N$412 VDD p l=2e-06 w=5e-06
M_MP347 N$14089 N$11347 N$412 VDD p l=2e-06 w=5e-06
M_MP346 N$324 N$14095 N$376 VDD p l=2e-06 w=5e-06
M_MP422 N$1652 N$1653 N$1655 VDD p l=2e-06 w=3e-06
M_MP421 N$1655 N$1653 VDD VDD p l=2e-06 w=3e-06
M_MP420 N$1655 N$11561 VDD VDD p l=2e-06 w=3e-06
M_MP444 N$1628 N$1636 N$1629 VDD p l=2e-06 w=3e-06
M_MP443 N$1629 N$11786 N$1630 VDD p l=2e-06 w=3e-06
M_MP419 N$13038 N$1662 VDD VDD p l=2e-06 w=3e-06
M_MP480 N$1674 N$13447 N$1593 VDD p l=2e-06 w=5e-06
M_MP479 N$1654 N$13243 N$1593 VDD p l=2e-06 w=5e-06
M_MP478 N$1654 N$13447 N$11816 VDD p l=2e-06 w=5e-06
M_MP483 N$1584 N$1589 VDD VDD p l=2e-06 w=6e-06
M_MP524 N$1549 N$1548 VDD VDD p l=2e-06 w=6e-06
M_MP764 N$11343 N$11342 VDD VDD p l=2e-06 w=6e-06
M_MP763 N$11344 N$11343 VDD VDD p l=2e-06 w=6e-06
M_MP762 N$11342 CK N$11344 VDD p l=2e-06 w=6e-06
M_MP761 N$11340 N$11339 N$11342 VDD p l=2e-06 w=6e-06
M_MP760 N$11340 N$11341 VDD VDD p l=2e-06 w=6e-06
M_MP539 N$14108 N$13857 VDD VDD p l=2e-06 w=6e-06
M_MP558 N$1521 CK N$1523 VDD p l=2e-06 w=6e-06
M_MP563 N$1517 CK SK0 VDD p l=2e-06 w=6e-06
M_MP536 N$1554 N$11083 VDD VDD p l=2e-06 w=6e-06
M_MP535 N$1540 CK N$1554 VDD p l=2e-06 w=6e-06
M_MP435 N$1638 N$1636 VDD VDD p l=2e-06 w=3e-06
M_MP434 N$1638 N$11786 VDD VDD p l=2e-06 w=3e-06
M_MP439 N$1633 N$1634 VDD VDD p l=2e-06 w=3e-06
M_MP470 N$1599 N$13243 N$1595 VDD p l=2e-06 w=5e-06
M_MP766 N$11345 N$11088 N$11108 VDD p l=2e-06 w=5e-06
M_MP521 N$13650 CK N$1552 VDD p l=2e-06 w=6e-06
M_MP413 N$1665 N$1654 VDD VDD p l=2e-06 w=3e-06
M_MP412 N$1665 N$11809 VDD VDD p l=2e-06 w=3e-06
M_MP504 N$1569 CK N$12429 VDD p l=2e-06 w=6e-06
M_MP472 N$13243 N$13447 VDD VDD p l=2e-06 w=5e-06
M_MP389 N$11780 CK VDD VDD p l=2e-06 w=5e-06
M_MP477 N$11561 N$13243 N$11816 VDD p l=2e-06 w=5e-06
M_MP476 N$11561 N$13447 N$11817 VDD p l=2e-06 w=5e-06
M_MP475 N$11786 N$13243 N$11817 VDD p l=2e-06 w=5e-06
M_MP488 N$1581 N$1583 VDD VDD p l=2e-06 w=6e-06
M_MP487 N$11571 N$1581 VDD VDD p l=2e-06 w=6e-06
M_MP507 N$1572 CK VDD VDD p l=2e-06 w=5e-06
M_MP506 N$12633 N$1569 VDD VDD p l=2e-06 w=6e-06
M_MP446 N$1627 N$1634 N$1630 VDD p l=2e-06 w=3e-06
M_MP445 N$1627 N$1650 N$1628 VDD p l=2e-06 w=3e-06
M_MP523 N$1548 N$1552 VDD VDD p l=2e-06 w=6e-06
M_MP522 N$1552 N$1551 N$1549 VDD p l=2e-06 w=6e-06
M_MP485 N$1585 N$1588 N$1583 VDD p l=2e-06 w=6e-06
M_MP469 N$13650 N$12835 N$1602 VDD p l=2e-06 w=6e-06
M_MP461 N$13039 N$1611 VDD VDD p l=2e-06 w=3e-06
M_MP433 N$13037 N$1644 VDD VDD p l=2e-06 w=3e-06
M_MP438 N$1634 N$11786 N$1635 VDD p l=2e-06 w=3e-06
M_MP437 N$1634 N$1650 N$1638 VDD p l=2e-06 w=3e-06
M_MP436 N$1635 N$1636 N$1638 VDD p l=2e-06 w=3e-06
M_MP94 N$94 N$90 VDD VDD p l=2e-06 w=3e-06
M_MP291 N$328 N$329 VDD VDD p l=2e-06 w=6e-06
M_MP344 N$317 N$14095 N$411 VDD p l=2e-06 w=5e-06
M_MP289 N$326 N$327 N$328 VDD p l=2e-06 w=6e-06
M_MP499 N$1595 CK N$1573 VDD p l=2e-06 w=6e-06
M_MP456 N$1614 N$1620 VDD VDD p l=2e-06 w=3e-06
M_MP455 N$1614 N$1599 VDD VDD p l=2e-06 w=3e-06
M_MP454 N$1614 N$1633 VDD VDD p l=2e-06 w=3e-06
M_MP453 N$13447 N$9715 VDD VDD p l=2e-06 w=3e-06
M_MP265 N$307 N$306 N$309 VDD p l=2e-06 w=6e-06
M_MP264 N$307 N$308 VDD VDD p l=2e-06 w=6e-06
M_MP263 N$308 N$305 VDD VDD p l=2e-06 w=6e-06
M_MP240 N$417 N$420 VDD VDD p l=2e-06 w=6e-06
M_MP429 N$1646 N$11561 N$1647 VDD p l=2e-06 w=3e-06
M_MP430 N$1645 N$1653 N$1646 VDD p l=2e-06 w=3e-06
M_MP591 SK3 N$1491 VDD VDD p l=2e-06 w=6e-06
M_MP590 N$1493 CK SK3 VDD p l=2e-06 w=6e-06
M_MP589 N$1495 N$1497 N$1493 VDD p l=2e-06 w=6e-06
M_MP562 N$1519 N$1522 N$1517 VDD p l=2e-06 w=6e-06
M_MP153 N$170 N$390 N$168 VDD p l=2e-06 w=3e-06
M_MP152 N$168 N$390 VDD VDD p l=2e-06 w=3e-06
M_MP275 N$316 CK N$317 VDD p l=2e-06 w=6e-06
M_MP274 N$314 N$313 N$316 VDD p l=2e-06 w=6e-06
M_MP273 N$314 N$315 VDD VDD p l=2e-06 w=6e-06
M_MP246 N$293 N$294 VDD VDD p l=2e-06 w=6e-06
M_MP217 N$183 N$14095 N$250 VDD p l=2e-06 w=5e-06
M_MP245 N$294 N$291 VDD VDD p l=2e-06 w=6e-06
M_MP244 N$291 N$292 N$293 VDD p l=2e-06 w=6e-06
M_MP288 N$258 CK N$326 VDD p l=2e-06 w=6e-06
M_MP298 N$333 N$334 N$335 VDD p l=2e-06 w=6e-06
M_MP87 N$87 0 VDD VDD p l=2e-06 w=3e-06
M_MP86 N$84 N$81 VDD VDD p l=2e-06 w=3e-06
M_MP460 N$1611 N$9715 N$1614 VDD p l=2e-06 w=3e-06
M_MP459 N$1611 N$1633 N$1612 VDD p l=2e-06 w=3e-06
M_MP458 N$1612 N$1620 N$1613 VDD p l=2e-06 w=3e-06
M_MP432 N$1644 N$1651 N$1647 VDD p l=2e-06 w=3e-06
M_MP431 N$1644 N$1668 N$1645 VDD p l=2e-06 w=3e-06
M_MP492 N$1577 N$1580 VDD VDD p l=2e-06 w=6e-06
M_MP491 N$1580 N$1579 N$1578 VDD p l=2e-06 w=6e-06
M_MP490 N$11816 CK N$1580 VDD p l=2e-06 w=6e-06
M_MP495 N$1576 CK N$11572 VDD p l=2e-06 w=6e-06
M_MP239 N$420 N$386 N$278 VDD p l=2e-06 w=6e-06
M_MP238 N$278 N$279 VDD VDD p l=2e-06 w=6e-06
M_MP258 N$384 N$304 VDD VDD p l=2e-06 w=6e-06
M_MP257 N$302 CK N$384 VDD p l=2e-06 w=6e-06
M_MP282 N$321 N$322 VDD VDD p l=2e-06 w=6e-06
M_MP501 N$1570 N$1573 VDD VDD p l=2e-06 w=6e-06
M_MP500 N$1573 N$1572 N$1571 VDD p l=2e-06 w=6e-06
M_MP532 N$1541 N$1545 VDD VDD p l=2e-06 w=6e-06
M_MP531 N$1545 N$1544 N$1542 VDD p l=2e-06 w=6e-06
M_MP503 N$1571 N$1572 N$1569 VDD p l=2e-06 w=6e-06
M_MP276 N$317 N$318 VDD VDD p l=2e-06 w=6e-06
M_MP561 N$1519 N$1518 VDD VDD p l=2e-06 w=6e-06
M_MP566 N$1522 CK VDD VDD p l=2e-06 w=5e-06
M_MP565 N$1515 N$1517 VDD VDD p l=2e-06 w=6e-06
M_MP564 SK0 N$1515 VDD VDD p l=2e-06 w=6e-06
M_MP410 N$1671 N$1654 N$1672 VDD p l=2e-06 w=3e-06
M_MP243 N$237 CK N$291 VDD p l=2e-06 w=6e-06
M_MP406 N$1675 N$1654 VDD VDD p l=2e-06 w=3e-06
M_MP262 N$305 N$306 N$307 VDD p l=2e-06 w=6e-06
M_MP261 N$246 CK N$305 VDD p l=2e-06 w=6e-06
M_MP411 N$1668 N$1671 VDD VDD p l=2e-06 w=3e-06
M_MP602 0 N$1557 N$1484 VDD p l=2e-06 w=5e-06
M_MP579 N$1503 N$1502 VDD VDD p l=2e-06 w=6e-06
M_MP486 N$1583 CK N$11571 VDD p l=2e-06 w=6e-06
M_MP577 N$1506 N$1505 N$1503 VDD p l=2e-06 w=6e-06
M_MP576 N$1504 CK N$1506 VDD p l=2e-06 w=6e-06
M_MP582 SK2 N$1499 VDD VDD p l=2e-06 w=6e-06
M_MP581 N$1501 CK SK2 VDD p l=2e-06 w=6e-06
M_MP580 N$1503 N$1505 N$1501 VDD p l=2e-06 w=6e-06
M_MP494 N$1578 N$1579 N$1576 VDD p l=2e-06 w=6e-06
M_MP260 N$299 CK VDD VDD p l=2e-06 w=5e-06
M_MP259 N$304 N$302 VDD VDD p l=2e-06 w=6e-06
M_MP498 N$1579 CK VDD VDD p l=2e-06 w=5e-06
M_MP497 N$1574 N$1576 VDD VDD p l=2e-06 w=6e-06
M_MP496 N$11572 N$1574 VDD VDD p l=2e-06 w=6e-06
M_MP585 N$1496 CK N$1498 VDD p l=2e-06 w=6e-06
M_MP618 N$1466 N$1465 VDD VDD p l=2e-06 w=3e-06
M_MP617 N$1466 B1 VDD VDD p l=2e-06 w=3e-06
M_MP623 N$1459 N$1477 VDD VDD p l=2e-06 w=3e-06
M_MP622 N$1462 N$1463 VDD VDD p l=2e-06 w=3e-06
M_MP594 N$11571 N$1489 N$1488 VDD p l=2e-06 w=5e-06
M_MP593 N$1497 CK VDD VDD p l=2e-06 w=5e-06
M_MP592 N$1491 N$1493 VDD VDD p l=2e-06 w=6e-06
M_MP597 N$11572 N$1489 N$1486 VDD p l=2e-06 w=5e-06
M_MP570 N$1511 N$1510 VDD VDD p l=2e-06 w=6e-06
M_MP569 N$1510 N$1514 VDD VDD p l=2e-06 w=6e-06
M_MP409 N$1671 N$11809 N$1675 VDD p l=2e-06 w=3e-06
M_MP408 N$1672 N$1673 N$1675 VDD p l=2e-06 w=3e-06
M_MP407 N$1675 N$1673 VDD VDD p l=2e-06 w=3e-06
M_MP573 SK1 N$1507 VDD VDD p l=2e-06 w=6e-06
M_MP572 N$1509 CK SK1 VDD p l=2e-06 w=6e-06
M_MP571 N$1511 N$1513 N$1509 VDD p l=2e-06 w=6e-06
M_MP635 N$1448 B2 N$1449 VDD p l=2e-06 w=3e-06
M_MP641 N$1442 N$1450 N$1443 VDD p l=2e-06 w=3e-06
M_MP640 N$1443 B2 N$1444 VDD p l=2e-06 w=3e-06
M_MP639 N$1444 N$1450 VDD VDD p l=2e-06 w=3e-06
M_MP638 N$1444 B2 VDD VDD p l=2e-06 w=3e-06
M_MP607 N$1479 B0 N$1480 VDD p l=2e-06 w=3e-06
M_MP606 N$1479 C N$1482 VDD p l=2e-06 w=3e-06
M_MP578 N$1502 N$1506 VDD VDD p l=2e-06 w=6e-06
M_MP610 N$1474 B0 VDD VDD p l=2e-06 w=3e-06
M_MP609 N$1474 C VDD VDD p l=2e-06 w=3e-06
M_MP608 N$1477 N$1479 VDD VDD p l=2e-06 w=3e-06
M_MP493 N$1578 N$1577 VDD VDD p l=2e-06 w=6e-06
M_MP583 N$1499 N$1501 VDD VDD p l=2e-06 w=6e-06
M_MP588 N$1495 N$1494 VDD VDD p l=2e-06 w=6e-06
M_MP587 N$1494 N$1498 VDD VDD p l=2e-06 w=6e-06
M_MP586 N$1498 N$1497 N$1495 VDD p l=2e-06 w=6e-06
M_MP620 N$1463 N$1477 N$1466 VDD p l=2e-06 w=3e-06
M_MP619 N$1464 N$1465 N$1466 VDD p l=2e-06 w=3e-06
M_MP657 N$1426 N$1433 N$1429 VDD p l=2e-06 w=3e-06
M_MP628 N$1456 N$1477 N$1457 VDD p l=2e-06 w=3e-06
M_MP627 N$1457 N$1465 N$1458 VDD p l=2e-06 w=3e-06
M_MP626 N$1458 B1 N$1459 VDD p l=2e-06 w=3e-06
M_MP625 N$1459 N$1465 VDD VDD p l=2e-06 w=3e-06
M_MP624 N$1459 B1 VDD VDD p l=2e-06 w=3e-06
M_MP596 N$1489 N$1557 VDD VDD p l=2e-06 w=5e-06
M_MP595 0 N$1557 N$1488 VDD p l=2e-06 w=5e-06
M_MP568 N$1514 N$1513 N$1511 VDD p l=2e-06 w=6e-06
M_MP567 N$1512 CK N$1514 VDD p l=2e-06 w=6e-06
M_MP599 N$12632 N$1489 N$1485 VDD p l=2e-06 w=5e-06
M_MP598 0 N$1557 N$1486 VDD p l=2e-06 w=5e-06
M_MP605 N$1480 N$1481 N$1482 VDD p l=2e-06 w=3e-06
M_MP604 N$1482 N$1481 VDD VDD p l=2e-06 w=3e-06
M_MP603 N$1482 B0 VDD VDD p l=2e-06 w=3e-06
M_MP667 N$1527 N$1557 N$1512 VDD p l=2e-06 w=5e-06
M_MP672 N$1467 N$1413 N$14097 VDD p l=2e-06 w=5e-06
M_MP637 N$1444 N$1462 VDD VDD p l=2e-06 w=3e-06
M_MP636 N$1447 N$1448 VDD VDD p l=2e-06 w=3e-06
M_MP611 N$1474 N$1481 VDD VDD p l=2e-06 w=3e-06
M_MP643 N$1441 N$1448 N$1444 VDD p l=2e-06 w=3e-06
M_MP642 N$1441 N$1462 N$1442 VDD p l=2e-06 w=3e-06
M_MP645 N$1436 B3 VDD VDD p l=2e-06 w=3e-06
M_MP615 N$1471 N$1479 N$1474 VDD p l=2e-06 w=3e-06
M_MP614 N$1471 C N$1472 VDD p l=2e-06 w=3e-06
M_MP613 N$1472 N$1481 N$1473 VDD p l=2e-06 w=3e-06
M_MP584 N$1505 CK VDD VDD p l=2e-06 w=5e-06
M_MP621 N$1463 B1 N$1464 VDD p l=2e-06 w=3e-06
M_MP650 CoutHK_SK N$1433 VDD VDD p l=2e-06 w=3e-06
M_MP684 N$1404 N$1403 VDD VDD p l=2e-06 w=6e-06
M_MP683 N$1403 N$1406 VDD VDD p l=2e-06 w=6e-06
M_MP682 N$1406 N$14098 N$1404 VDD p l=2e-06 w=6e-06
M_MP656 N$1426 N$1447 N$1427 VDD p l=2e-06 w=3e-06
M_MP655 N$1427 N$1435 N$1428 VDD p l=2e-06 w=3e-06
M_MP654 N$1428 B3 N$1429 VDD p l=2e-06 w=3e-06
M_MP629 N$1456 N$1463 N$1459 VDD p l=2e-06 w=3e-06
M_MP658 N$1422 N$1426 VDD VDD p l=2e-06 w=3e-06
M_MP661 N$1435 N$1484 VDD VDD p l=2e-06 w=3e-06
M_MP601 N$12429 N$1489 N$1484 VDD p l=2e-06 w=5e-06
M_MP600 0 N$1557 N$1485 VDD p l=2e-06 w=5e-06
M_MP632 N$1451 N$1450 VDD VDD p l=2e-06 w=3e-06
M_MP631 N$1451 B2 VDD VDD p l=2e-06 w=3e-06
M_MP630 N$1452 N$1456 VDD VDD p l=2e-06 w=3e-06
M_MP668 N$1485 N$1416 N$1504 VDD p l=2e-06 w=5e-06
M_MP699 N$1409 CK N$1394 VDD p l=2e-06 w=6e-06
M_MP698 N$1399 CK VDD VDD p l=2e-06 w=5e-06
M_MP671 N$1525 N$1557 N$1496 VDD p l=2e-06 w=5e-06
M_MP340 N$384 N$14095 N$410 VDD p l=2e-06 w=5e-06
M_MP339 N$14085 N$11347 N$410 VDD p l=2e-06 w=5e-06
M_MP358 P2 N$409 N$387 VDD p l=2e-06 w=5e-06
M_MP355 N$409 N$14096 VDD VDD p l=2e-06 w=5e-06
M_MP678 0 N$1557 N$1409 VDD p l=2e-06 w=5e-06
M_MP612 N$1473 B0 N$1474 VDD p l=2e-06 w=3e-06
M_MP616 N$1467 N$1471 VDD VDD p l=2e-06 w=3e-06
M_MP649 N$1433 B3 N$1434 VDD p l=2e-06 w=3e-06
M_MP648 N$1433 N$1447 N$1436 VDD p l=2e-06 w=3e-06
M_MP647 N$1434 N$1435 N$1436 VDD p l=2e-06 w=3e-06
M_MP646 N$1436 N$1435 VDD VDD p l=2e-06 w=3e-06
M_MP652 N$1429 B3 VDD VDD p l=2e-06 w=3e-06
M_MP651 N$1429 N$1447 VDD VDD p l=2e-06 w=3e-06
M_MP679 N$1422 N$1413 N$1408 VDD p l=2e-06 w=5e-06
M_MP716 N$1387 CK VDD VDD p l=2e-06 w=5e-06
M_MP715 N$1383 N$1384 VDD VDD p l=2e-06 w=6e-06
M_MP714 N$14092 N$1383 VDD VDD p l=2e-06 w=6e-06
M_MP688 N$1401 N$1402 VDD VDD p l=2e-06 w=6e-06
M_MP687 N$14046 N$1401 VDD VDD p l=2e-06 w=6e-06
M_MP653 N$1429 N$1435 VDD VDD p l=2e-06 w=3e-06
M_MP399 N$11799 N$1674 VDD VDD p l=2e-06 w=3e-06
M_MP398 N$11799 C VDD VDD p l=2e-06 w=3e-06
M_MP397 N$11809 N$11796 VDD VDD p l=2e-06 w=3e-06
M_MP634 N$1448 N$1462 N$1451 VDD p l=2e-06 w=3e-06
M_MP633 N$1449 N$1450 N$1451 VDD p l=2e-06 w=3e-06
M_MP665 N$1416 N$1557 VDD VDD p l=2e-06 w=5e-06
M_MP664 N$1529 N$1557 N$1521 VDD p l=2e-06 w=5e-06
M_MP669 N$1526 N$1557 N$1504 VDD p l=2e-06 w=5e-06
M_MP556 N$12632 N$1530 N$1525 VDD p l=2e-06 w=5e-06
M_MP555 0 N$14108 N$1526 VDD p l=2e-06 w=5e-06
M_MP560 N$1518 N$1523 VDD VDD p l=2e-06 w=6e-06
M_MP559 N$1523 N$1522 N$1519 VDD p l=2e-06 w=6e-06
M_MP489 N$1588 CK VDD VDD p l=2e-06 w=5e-06
M_MP778 N$13885 N$14085 VDD VDD p l=2e-06 w=3e-06
M_MP777 OUT0 N$13879 VDD VDD p l=2e-06 w=3e-06
M_MP575 N$1513 CK VDD VDD p l=2e-06 w=5e-06
M_MP677 N$1437 N$1413 N$1409 VDD p l=2e-06 w=5e-06
M_MP676 0 N$1557 N$1410 VDD p l=2e-06 w=5e-06
M_MP712 N$1386 N$1387 N$1384 VDD p l=2e-06 w=6e-06
M_MP711 N$1386 N$1385 VDD VDD p l=2e-06 w=6e-06
M_MP511 N$13870 N$14084 N$13869 VDD p l=2e-06 w=3e-06
M_MP510 N$13870 0 N$13868 VDD p l=2e-06 w=3e-06
M_MP509 N$13869 N$13996 N$13868 VDD p l=2e-06 w=3e-06
M_MP508 N$13868 N$13996 VDD VDD p l=2e-06 w=3e-06
M_MP474 N$13868 N$14084 VDD VDD p l=2e-06 w=3e-06
M_MP400 N$11799 N$11794 VDD VDD p l=2e-06 w=3e-06
M_MP794 N$13902 N$14001 N$13901 VDD p l=2e-06 w=3e-06
M_MP793 N$13901 N$14001 VDD VDD p l=2e-06 w=3e-06
M_MP792 N$13901 N$14086 VDD VDD p l=2e-06 w=3e-06
M_MP791 OUT1 N$13895 VDD VDD p l=2e-06 w=3e-06
M_MP396 N$11796 N$1674 N$11795 VDD p l=2e-06 w=3e-06
M_MP395 N$11796 C N$11793 VDD p l=2e-06 w=3e-06
M_MP235 N$421 N$385 N$274 VDD p l=2e-06 w=6e-06
M_MP234 N$274 N$275 VDD VDD p l=2e-06 w=6e-06
M_MP553 0 N$14108 N$1527 VDD p l=2e-06 w=5e-06
M_MP552 N$11571 N$1530 N$1527 VDD p l=2e-06 w=5e-06
M_MP557 0 N$14108 N$1525 VDD p l=2e-06 w=5e-06
M_MP783 N$13889 N$13887 VDD VDD p l=2e-06 w=3e-06
M_MP782 N$13887 N$14085 N$13886 VDD p l=2e-06 w=3e-06
M_MP781 N$13887 N$13873 N$13885 VDD p l=2e-06 w=3e-06
M_MP780 N$13886 N$14000 N$13885 VDD p l=2e-06 w=3e-06
M_MP779 N$13885 N$14000 VDD VDD p l=2e-06 w=3e-06
M_MP810 N$13919 N$14087 N$13918 VDD p l=2e-06 w=3e-06
M_MP809 N$13919 N$13905 N$13917 VDD p l=2e-06 w=3e-06
M_MP808 N$13918 N$14002 N$13917 VDD p l=2e-06 w=3e-06
M_MP807 N$13917 N$14002 VDD VDD p l=2e-06 w=3e-06
M_MP806 N$13917 N$14087 VDD VDD p l=2e-06 w=3e-06
M_MP554 N$11572 N$1530 N$1526 VDD p l=2e-06 w=5e-06
M_MP774 N$13878 N$13996 N$13877 VDD p l=2e-06 w=3e-06
M_MP516 N$13877 N$14084 N$13876 VDD p l=2e-06 w=3e-06
M_MP515 N$13876 N$13996 VDD VDD p l=2e-06 w=3e-06
M_MP514 N$13876 N$14084 VDD VDD p l=2e-06 w=3e-06
M_MP513 N$13876 0 VDD VDD p l=2e-06 w=3e-06
M_MP512 N$13873 N$13870 VDD VDD p l=2e-06 w=3e-06
M_MP799 N$13908 N$14086 VDD VDD p l=2e-06 w=3e-06
M_MP798 N$13908 N$13889 VDD VDD p l=2e-06 w=3e-06
M_MP797 N$13905 N$13903 VDD VDD p l=2e-06 w=3e-06
M_MP796 N$13903 N$14086 N$13902 VDD p l=2e-06 w=3e-06
M_MP795 N$13903 N$13889 N$13901 VDD p l=2e-06 w=3e-06
M_MP824 N$13935 N$14088 N$13934 VDD p l=2e-06 w=3e-06
M_MP823 N$13935 N$13921 N$13933 VDD p l=2e-06 w=3e-06
M_MP822 N$13934 N$14003 N$13933 VDD p l=2e-06 w=3e-06
M_MP821 N$13933 N$14003 VDD VDD p l=2e-06 w=3e-06
M_MP820 N$13933 N$14088 VDD VDD p l=2e-06 w=3e-06
M_MP394 N$11795 N$11794 N$11793 VDD p l=2e-06 w=3e-06
M_MP393 N$11793 N$11794 VDD VDD p l=2e-06 w=3e-06
M_MP392 N$11793 N$1674 VDD VDD p l=2e-06 w=3e-06
M_MP790 N$13895 N$13887 N$13892 VDD p l=2e-06 w=3e-06
M_MP789 N$13895 N$13873 N$13894 VDD p l=2e-06 w=3e-06
M_MP788 N$13894 N$14000 N$13893 VDD p l=2e-06 w=3e-06
M_MP787 N$13893 N$14085 N$13892 VDD p l=2e-06 w=3e-06
M_MP786 N$13892 N$14000 VDD VDD p l=2e-06 w=3e-06
M_MP785 N$13892 N$14085 VDD VDD p l=2e-06 w=3e-06
M_MP784 N$13892 N$13873 VDD VDD p l=2e-06 w=3e-06
M_MP815 N$13925 N$14087 N$13924 VDD p l=2e-06 w=3e-06
M_MP814 N$13924 N$14002 VDD VDD p l=2e-06 w=3e-06
M_MP813 N$13924 N$14087 VDD VDD p l=2e-06 w=3e-06
M_MP812 N$13924 N$13905 VDD VDD p l=2e-06 w=3e-06
M_MP811 N$13921 N$13919 VDD VDD p l=2e-06 w=3e-06
M_MP838 N$13951 N$14089 N$13950 VDD p l=2e-06 w=3e-06
M_MP837 N$13951 N$13937 N$13949 VDD p l=2e-06 w=3e-06
M_MP836 N$13950 N$14004 N$13949 VDD p l=2e-06 w=3e-06
M_MP835 N$13949 N$14004 VDD VDD p l=2e-06 w=3e-06
M_MP805 OUT2 N$13911 VDD VDD p l=2e-06 w=3e-06
M_MP776 N$13879 N$13870 N$13876 VDD p l=2e-06 w=3e-06
M_MP775 N$13879 0 N$13878 VDD p l=2e-06 w=3e-06
M_MP804 N$13911 N$13903 N$13908 VDD p l=2e-06 w=3e-06
M_MP803 N$13911 N$13889 N$13910 VDD p l=2e-06 w=3e-06
M_MP802 N$13910 N$14001 N$13909 VDD p l=2e-06 w=3e-06
M_MP801 N$13909 N$14086 N$13908 VDD p l=2e-06 w=3e-06
M_MP800 N$13908 N$14001 VDD VDD p l=2e-06 w=3e-06
M_MP831 N$13943 N$13921 N$13942 VDD p l=2e-06 w=3e-06
M_MP830 N$13942 N$14003 N$13941 VDD p l=2e-06 w=3e-06
M_MP829 N$13941 N$14088 N$13940 VDD p l=2e-06 w=3e-06
M_MP828 N$13940 N$14003 VDD VDD p l=2e-06 w=3e-06
M_MP827 N$13940 N$14088 VDD VDD p l=2e-06 w=3e-06
M_MP826 N$13940 N$13921 VDD VDD p l=2e-06 w=3e-06
M_MP825 N$13937 N$13935 VDD VDD p l=2e-06 w=3e-06
M_MP852 N$13967 N$14090 N$13966 VDD p l=2e-06 w=3e-06
M_MP851 N$13967 N$13953 N$13965 VDD p l=2e-06 w=3e-06
M_MP819 OUT3 N$13927 VDD VDD p l=2e-06 w=3e-06
M_MP818 N$13927 N$13919 N$13924 VDD p l=2e-06 w=3e-06
M_MP817 N$13927 N$13905 N$13926 VDD p l=2e-06 w=3e-06
M_MP816 N$13926 N$14002 N$13925 VDD p l=2e-06 w=3e-06
M_MP846 N$13959 N$13951 N$13956 VDD p l=2e-06 w=3e-06
M_MP845 N$13959 N$13937 N$13958 VDD p l=2e-06 w=3e-06
M_MP844 N$13958 N$14004 N$13957 VDD p l=2e-06 w=3e-06
M_MP843 N$13957 N$14089 N$13956 VDD p l=2e-06 w=3e-06
M_MP842 N$13956 N$14004 VDD VDD p l=2e-06 w=3e-06
M_MP841 N$13956 N$14089 VDD VDD p l=2e-06 w=3e-06
M_MP840 N$13956 N$13937 VDD VDD p l=2e-06 w=3e-06
M_MP839 N$13953 N$13951 VDD VDD p l=2e-06 w=3e-06
M_MP868 N$13988 N$13969 VDD VDD p l=2e-06 w=3e-06
M_MP867 CARRY_OUT N$13983 VDD VDD p l=2e-06 w=3e-06
M_MP834 N$13949 N$14089 VDD VDD p l=2e-06 w=3e-06
M_MP832 N$13943 N$13935 N$13940 VDD p l=2e-06 w=3e-06
M_MP860 N$13975 N$13967 N$13972 VDD p l=2e-06 w=3e-06
M_MP859 N$13975 N$13953 N$13974 VDD p l=2e-06 w=3e-06
M_MP858 N$13974 N$14005 N$13973 VDD p l=2e-06 w=3e-06
M_MP857 N$13973 N$14090 N$13972 VDD p l=2e-06 w=3e-06
M_MP856 N$13972 N$14005 VDD VDD p l=2e-06 w=3e-06
M_MP855 N$13972 N$14090 VDD VDD p l=2e-06 w=3e-06
M_MP854 N$13972 N$13953 VDD VDD p l=2e-06 w=3e-06
M_MP853 N$13969 N$13967 VDD VDD p l=2e-06 w=3e-06
M_MP930 N$14014 SK3 N$14005 VDD p l=2e-06 w=5e-06
M_MP929 N$14006 SK3 VDD VDD p l=2e-06 w=5e-06
M_MP934 N$14012 SK3 N$14003 VDD p l=2e-06 w=5e-06
M_MP933 N$14010 N$14006 N$14004 VDD p l=2e-06 w=5e-06
M_MP900 N$14031 SK1 N$14021 VDD p l=2e-06 w=5e-06
M_MP847 OUT5 N$13959 VDD VDD p l=2e-06 w=3e-06
M_MP874 N$13991 N$13983 N$13988 VDD p l=2e-06 w=3e-06
M_MP873 N$13991 N$13969 N$13990 VDD p l=2e-06 w=3e-06
M_MP872 N$13990 N$14007 N$13989 VDD p l=2e-06 w=3e-06
M_MP871 N$13989 N$14091 N$13988 VDD p l=2e-06 w=3e-06
M_MP870 N$13988 N$14007 VDD VDD p l=2e-06 w=3e-06
M_MP869 N$13988 N$14091 VDD VDD p l=2e-06 w=3e-06
M_MP947 N$13997 N$11347 N$13998 VDD p l=2e-06 w=5e-06
M_MP946 N$13998 N$11083 VDD VDD p l=2e-06 w=5e-06
M_MP945 N$13999 N$14108 N$14040 VDD p l=2e-06 w=5e-06
M_MP948 N$13999 N$13997 VDD VDD p l=2e-06 w=5e-06
M_MP916 N$14020 N$14015 N$14013 VDD p l=2e-06 w=5e-06
M_MP833 OUT4 N$13943 VDD VDD p l=2e-06 w=3e-06
M_MP861 OUT6 N$13975 VDD VDD p l=2e-06 w=3e-06
M_MP923 N$14018 SK2 N$14009 VDD p l=2e-06 w=5e-06
M_MP922 N$14017 N$14015 N$14010 VDD p l=2e-06 w=5e-06
M_MP928 N$14012 N$14006 N$14007 VDD p l=2e-06 w=5e-06
M_MP927 N$14016 SK3 N$14007 VDD p l=2e-06 w=5e-06
M_MP926 0 N$14015 N$14008 VDD p l=2e-06 w=5e-06
M_MP925 N$14017 SK2 N$14008 VDD p l=2e-06 w=5e-06
M_MP931 N$14011 N$14006 N$14005 VDD p l=2e-06 w=5e-06
M_MP222 N$200 N$265 N$258 VDD p l=2e-06 w=5e-06
M_MP418 N$1662 N$1671 N$1665 VDD p l=2e-06 w=3e-06
M_MP417 N$1662 N$11809 N$1663 VDD p l=2e-06 w=3e-06
M_MP416 N$1663 N$1673 N$1664 VDD p l=2e-06 w=3e-06
M_MP415 N$1664 N$1654 N$1665 VDD p l=2e-06 w=3e-06
M_MP299 N$336 N$333 VDD VDD p l=2e-06 w=6e-06
M_MP266 N$309 CK N$310 VDD p l=2e-06 w=6e-06
M_MP232 N$112 N$14095 N$271 VDD p l=2e-06 w=5e-06
M_MP905 N$14028 N$14024 N$14019 VDD p l=2e-06 w=5e-06
M_MP904 N$14029 SK1 N$14019 VDD p l=2e-06 w=5e-06
M_MP903 N$14029 N$14024 N$14020 VDD p l=2e-06 w=5e-06
M_MP908 N$14027 SK1 N$14017 VDD p l=2e-06 w=5e-06
M_MP939 0 N$14006 N$14001 VDD p l=2e-06 w=5e-06
M_MP938 N$14010 SK3 N$14001 VDD p l=2e-06 w=5e-06
M_MP944 N$11083 N$13857 N$14040 VDD p l=2e-06 w=5e-06
M_MP943 0 N$14006 N$13996 VDD p l=2e-06 w=5e-06
M_MP942 N$14008 SK3 N$13996 VDD p l=2e-06 w=5e-06
M_MP941 0 N$14006 N$14000 VDD p l=2e-06 w=5e-06
M_MP197 N$222 N$14081 N$221 VDD p l=2e-06 w=3e-06
M_MP151 N$168 N$14078 VDD VDD p l=2e-06 w=3e-06
M_MP131 N$141 N$388 VDD VDD p l=2e-06 w=3e-06
M_MP122 N$130 N$126 VDD VDD p l=2e-06 w=3e-06
M_MP921 N$14019 SK2 N$14010 VDD p l=2e-06 w=5e-06
M_MP920 N$14018 N$14015 N$14011 VDD p l=2e-06 w=5e-06
M_MP919 N$14020 SK2 N$14011 VDD p l=2e-06 w=5e-06
M_MP924 0 N$14015 N$14009 VDD p l=2e-06 w=5e-06
M_MP130 N$141 0 VDD VDD p l=2e-06 w=3e-06
M_MP129 N$141 N$120 VDD VDD p l=2e-06 w=3e-06
M_MP128 N$138 N$136 VDD VDD p l=2e-06 w=3e-06
M_MP172 N$193 N$14079 VDD VDD p l=2e-06 w=3e-06
M_MP201 N$227 N$395 VDD VDD p l=2e-06 w=3e-06
M_MP200 N$227 N$14081 VDD VDD p l=2e-06 w=3e-06
M_MP199 N$227 N$207 VDD VDD p l=2e-06 w=3e-06
M_MP198 Cout N$222 VDD VDD p l=2e-06 w=3e-06
M_MP223 N$217 N$14095 N$258 VDD p l=2e-06 w=5e-06
M_MP211 N$148 N$14095 N$242 VDD p l=2e-06 w=5e-06
M_MP210 N$130 N$265 N$242 VDD p l=2e-06 w=5e-06
M_MP168 N$188 N$173 N$185 VDD p l=2e-06 w=3e-06
M_MP167 N$187 N$392 N$185 VDD p l=2e-06 w=3e-06
M_MP108 N$112 N$108 VDD VDD p l=2e-06 w=3e-06
M_MP231 N$94 N$265 N$271 VDD p l=2e-06 w=5e-06
M_MP302 N$337 CK N$338 VDD p l=2e-06 w=6e-06
M_MP303 N$338 N$339 VDD VDD p l=2e-06 w=6e-06
M_MP206 N$1179 N$230 VDD VDD p l=2e-06 w=3e-06
M_MP237 N$275 N$386 VDD VDD p l=2e-06 w=6e-06
M_MP236 N$419 N$421 VDD VDD p l=2e-06 w=6e-06
M_MP256 N$300 N$299 N$302 VDD p l=2e-06 w=6e-06
M_MP185 N$210 N$190 VDD VDD p l=2e-06 w=3e-06
M_MP184 N$207 N$205 VDD VDD p l=2e-06 w=3e-06
M_MP99 N$100 0 N$99 VDD p l=2e-06 w=3e-06
M_MP12 N$15 N$17 VDD VDD p l=2e-06 w=6e-06
M_MP93 N$90 N$81 N$87 VDD p l=2e-06 w=3e-06
M_MP121 N$126 N$118 N$123 VDD p l=2e-06 w=3e-06
M_MP120 N$126 N$102 N$125 VDD p l=2e-06 w=3e-06
M_MP119 N$125 N$387 N$124 VDD p l=2e-06 w=3e-06
M_MP118 N$124 0 N$123 VDD p l=2e-06 w=3e-06
M_MP117 N$123 N$387 VDD VDD p l=2e-06 w=3e-06
M_MP546 N$11572 RST N$11561 VDD p l=2e-06 w=5e-06
M_MP545 0 N$11813 N$11561 VDD p l=2e-06 w=5e-06
M_MP544 N$11571 RST N$1654 VDD p l=2e-06 w=5e-06
M_MP543 0 N$11813 N$1654 VDD p l=2e-06 w=5e-06
M_MP377 N$11790 CK N$14107 VDD p l=2e-06 w=6e-06
M_MP181 N$204 N$394 N$202 VDD p l=2e-06 w=3e-06
M_MP136 N$148 N$144 VDD VDD p l=2e-06 w=3e-06
M_MP290 N$329 N$326 VDD VDD p l=2e-06 w=6e-06
M_MP316 N$361 N$11347 OUT8 VDD p l=2e-06 w=5e-06
M_MP309 N$342 N$343 VDD VDD p l=2e-06 w=6e-06
M_MP308 N$343 N$340 VDD VDD p l=2e-06 w=6e-06
M_MP307 N$340 N$341 N$342 VDD p l=2e-06 w=6e-06
M_MP306 N$266 CK N$340 VDD p l=2e-06 w=6e-06
M_MP101 N$105 N$84 VDD VDD p l=2e-06 w=3e-06
M_MP100 N$102 N$100 VDD VDD p l=2e-06 w=3e-06
M_MP156 N$173 N$171 VDD VDD p l=2e-06 w=3e-06
M_MP320 0 N$348 N$14085 VDD p l=2e-06 w=5e-06
M_MP329 0 N$348 N$14089 VDD p l=2e-06 w=5e-06
M_MP248 N$295 CK N$296 VDD p l=2e-06 w=6e-06
M_MP247 N$293 N$292 N$295 VDD p l=2e-06 w=6e-06
M_MP280 N$319 N$320 N$321 VDD p l=2e-06 w=6e-06
M_MP216 N$166 N$265 N$250 VDD p l=2e-06 w=5e-06
M_MP692 N$1397 N$1400 VDD VDD p l=2e-06 w=6e-06
M_MP109 N$114 0 VDD VDD p l=2e-06 w=3e-06
M_MP233 N$265 N$14095 VDD VDD p l=2e-06 w=5e-06
M_MP110 N$114 N$387 VDD VDD p l=2e-06 w=3e-06
M_MP208 N$130 N$14095 N$237 VDD p l=2e-06 w=5e-06
M_MP375 N$11783 N$11782 VDD VDD p l=2e-06 w=6e-06
M_MP374 N$11782 N$11784 VDD VDD p l=2e-06 w=6e-06
M_MP373 N$11784 N$11789 N$11783 VDD p l=2e-06 w=6e-06
M_MP372 N$11570 CK N$11784 VDD p l=2e-06 w=6e-06
M_MP64 N$286 N$287 VDD VDD p l=2e-06 w=6e-06
M_MP63 N$287 N$282 VDD VDD p l=2e-06 w=6e-06
M_MP192 N$217 N$213 VDD VDD p l=2e-06 w=3e-06
M_MP177 N$196 N$188 N$193 VDD p l=2e-06 w=3e-06
M_MP287 N$320 CK VDD VDD p l=2e-06 w=5e-06
M_MP214 N$166 N$14095 N$246 VDD p l=2e-06 w=5e-06
M_MP92 N$90 0 N$89 VDD p l=2e-06 w=3e-06
M_MP91 N$89 N$385 N$88 VDD p l=2e-06 w=3e-06
M_MP90 N$88 0 N$87 VDD p l=2e-06 w=3e-06
M_MP89 N$87 N$385 VDD VDD p l=2e-06 w=3e-06
M_MP88 N$87 0 VDD VDD p l=2e-06 w=3e-06
M_MP116 N$123 0 VDD VDD p l=2e-06 w=3e-06
M_MP115 N$123 N$102 VDD VDD p l=2e-06 w=3e-06
M_MP114 N$120 N$118 VDD VDD p l=2e-06 w=3e-06
M_MP142 N$156 N$154 VDD VDD p l=2e-06 w=3e-06
M_MP171 N$193 N$173 VDD VDD p l=2e-06 w=3e-06
M_MP170 N$190 N$188 VDD VDD p l=2e-06 w=3e-06
M_MP277 N$318 N$316 VDD VDD p l=2e-06 w=6e-06
M_MP250 N$297 N$295 VDD VDD p l=2e-06 w=6e-06
M_MP249 N$296 N$297 VDD VDD p l=2e-06 w=6e-06
M_MP331 0 N$348 N$14090 VDD p l=2e-06 w=5e-06
M_MP547 0 N$11813 N$11786 VDD p l=2e-06 w=5e-06
M_MP527 N$1558 N$1546 VDD VDD p l=2e-06 w=6e-06
M_MP281 N$322 N$319 VDD VDD p l=2e-06 w=6e-06
M_MP242 N$283 CK VDD VDD p l=2e-06 w=5e-06
M_MP68 N$290 N$288 VDD VDD p l=2e-06 w=6e-06
M_MP304 N$339 N$337 VDD VDD p l=2e-06 w=6e-06
M_MP278 N$313 CK VDD VDD p l=2e-06 w=5e-06
M_MP283 N$321 N$320 N$323 VDD p l=2e-06 w=6e-06
M_MP220 N$200 N$14095 N$254 VDD p l=2e-06 w=5e-06
M_MP219 N$183 N$265 N$254 VDD p l=2e-06 w=5e-06
M_MP279 N$254 CK N$319 VDD p l=2e-06 w=6e-06
M_MP352 N$345 N$14095 N$396 VDD p l=2e-06 w=5e-06
M_MP83 N$80 N$385 N$77 VDD p l=2e-06 w=3e-06
M_MP226 N$1179 N$14095 N$262 VDD p l=2e-06 w=5e-06
M_MP272 N$315 N$312 VDD VDD p l=2e-06 w=6e-06
M_MP163 N$179 N$171 N$176 VDD p l=2e-06 w=3e-06
M_MP162 N$179 N$156 N$178 VDD p l=2e-06 w=3e-06
M_MP169 N$188 N$14079 N$187 VDD p l=2e-06 w=3e-06
M_MP138 N$150 N$389 VDD VDD p l=2e-06 w=3e-06
M_MP137 N$150 0 VDD VDD p l=2e-06 w=3e-06
M_MP319 N$296 N$11347 N$14084 VDD p l=2e-06 w=5e-06
M_MP318 0 N$348 N$14084 VDD p l=2e-06 w=5e-06
M_MP317 N$348 N$11347 VDD VDD p l=2e-06 w=5e-06
M_MP769 N$11802 N$11796 N$11799 VDD p l=2e-06 w=3e-06
M_MP768 N$11802 C N$11801 VDD p l=2e-06 w=3e-06
M_MP402 N$11801 N$11794 N$11800 VDD p l=2e-06 w=3e-06
M_MP401 N$11800 N$1674 N$11799 VDD p l=2e-06 w=3e-06
M_MP452 N$9715 N$1599 N$1619 VDD p l=2e-06 w=3e-06
M_MP451 N$9715 N$1633 N$1622 VDD p l=2e-06 w=3e-06
M_MP457 N$1613 N$1599 N$1614 VDD p l=2e-06 w=3e-06
M_MP351 N$14091 N$11347 N$396 VDD p l=2e-06 w=5e-06
M_MP731 N$11324 CK N$11099 VDD p l=2e-06 w=6e-06
M_MP732 N$11099 N$11325 VDD VDD p l=2e-06 w=6e-06
M_MP721 N$11316 N$11315 N$11318 VDD p l=2e-06 w=6e-06
M_MP720 N$11316 N$11317 VDD VDD p l=2e-06 w=6e-06
M_MP719 N$11317 N$11314 VDD VDD p l=2e-06 w=6e-06
M_MP718 N$11314 N$11315 N$11316 VDD p l=2e-06 w=6e-06
M_MP717 N$382 CK N$11314 VDD p l=2e-06 w=6e-06
M_MP752 N$11334 N$11333 N$11336 VDD p l=2e-06 w=6e-06
M_MP442 N$1630 N$1636 VDD VDD p l=2e-06 w=3e-06
M_MP441 N$1630 N$11786 VDD VDD p l=2e-06 w=3e-06
M_MP440 N$1630 N$1650 VDD VDD p l=2e-06 w=3e-06
M_MP537 N$11083 N$1540 VDD VDD p l=2e-06 w=6e-06
M_MP534 N$1542 N$1544 N$1540 VDD p l=2e-06 w=6e-06
M_MP888 0 N$14037 N$14029 VDD p l=2e-06 w=5e-06
M_MP896 N$14035 SK1 N$14023 VDD p l=2e-06 w=5e-06
M_MP525 N$1549 N$1551 N$1547 VDD p l=2e-06 w=6e-06
M_MP530 N$13447 CK N$1545 VDD p l=2e-06 w=6e-06
M_MP529 N$1551 CK VDD VDD p l=2e-06 w=6e-06
M_MP528 N$1546 N$1547 VDD VDD p l=2e-06 w=6e-06
M_MP533 N$1542 N$1541 VDD VDD p l=2e-06 w=6e-06
M_MP473 N$13651 N$13039 VDD VDD p l=2e-06 w=5e-06
M_MP526 N$1547 CK N$1558 VDD p l=2e-06 w=6e-06
M_MP548 N$12632 RST N$11786 VDD p l=2e-06 w=5e-06
M_MP482 N$1589 N$1588 N$1585 VDD p l=2e-06 w=6e-06
M_MP481 N$1593 CK N$1589 VDD p l=2e-06 w=6e-06
M_MP877 0 N$14037 N$14039 VDD p l=2e-06 w=5e-06
M_MP876 0 N$14040 N$14039 VDD p l=2e-06 w=5e-06
M_MP906 N$14028 SK1 N$14018 VDD p l=2e-06 w=5e-06
M_MP912 N$14015 SK2 VDD VDD p l=2e-06 w=5e-06
M_MP911 N$14022 N$14015 N$14016 VDD p l=2e-06 w=5e-06
M_MP464 N$1620 0 VDD VDD p l=2e-06 w=3e-06
M_MP463 N$1653 B2 VDD VDD p l=2e-06 w=3e-06
M_MP462 N$1673 B1 VDD VDD p l=2e-06 w=3e-06
M_MP484 N$1585 N$1584 VDD VDD p l=2e-06 w=6e-06
M_MP468 N$1602 N$13037 N$1603 VDD p l=2e-06 w=6e-06
M_MP467 N$1603 N$13038 N$1604 VDD p l=2e-06 w=6e-06
M_MP466 N$1604 N$11810 N$13651 VDD p l=2e-06 w=6e-06
M_MP465 N$1636 B3 VDD VDD p l=2e-06 w=3e-06
M_MP471 N$11786 N$13447 N$1595 VDD p l=2e-06 w=5e-06
M_MP426 N$1647 N$1668 VDD VDD p l=2e-06 w=3e-06
M_MP425 N$1650 N$1651 VDD VDD p l=2e-06 w=3e-06
M_MP541 N$14107 RST N$1674 VDD p l=2e-06 w=5e-06
M_MP540 A5 N$11813 N$1674 VDD p l=2e-06 w=5e-06
M_MP414 N$1665 N$1673 VDD VDD p l=2e-06 w=3e-06
M_MP907 N$14027 N$14024 N$14018 VDD p l=2e-06 w=5e-06
M_MP890 0 N$14037 N$14028 VDD p l=2e-06 w=5e-06
M_MP889 P2 N$14040 N$14028 VDD p l=2e-06 w=5e-06
M_MP381 N$11817 CK N$11781 VDD p l=2e-06 w=6e-06
M_MP380 N$11789 CK VDD VDD p l=2e-06 w=5e-06
M_MP895 N$14024 SK1 VDD VDD p l=2e-06 w=5e-06
M_MP894 N$14035 N$14024 N$14025 VDD p l=2e-06 w=5e-06
M_MP899 N$14031 N$14024 N$14022 VDD p l=2e-06 w=5e-06
M_MP898 N$14033 SK1 N$14022 VDD p l=2e-06 w=5e-06
M_MP897 N$14033 N$14024 N$14023 VDD p l=2e-06 w=5e-06
M_MP902 N$14030 SK1 N$14020 VDD p l=2e-06 w=5e-06
M_MP901 N$14030 N$14024 N$14021 VDD p l=2e-06 w=5e-06
M_MP866 N$13983 N$14091 N$13982 VDD p l=2e-06 w=3e-06
M_MP865 N$13983 N$13969 N$13981 VDD p l=2e-06 w=3e-06
M_MP864 N$13982 N$14007 N$13981 VDD p l=2e-06 w=3e-06
M_MP863 N$13981 N$14007 VDD VDD p l=2e-06 w=3e-06
M_MP862 N$13981 N$14091 VDD VDD p l=2e-06 w=3e-06
M_MP878 N$14037 N$14040 VDD VDD p l=2e-06 w=5e-06
M_MP940 N$14009 SK3 N$14000 VDD p l=2e-06 w=5e-06
M_MP743 N$11327 CK VDD VDD p l=2e-06 w=5e-06
M_MP753 N$11336 CK N$382 VDD p l=2e-06 w=6e-06
M_MP910 N$14025 SK2 N$14016 VDD p l=2e-06 w=5e-06
M_MP909 0 N$14024 N$14017 VDD p l=2e-06 w=5e-06
M_MP915 N$14022 SK2 N$14013 VDD p l=2e-06 w=5e-06
M_MP914 N$14021 N$14015 N$14014 VDD p l=2e-06 w=5e-06
M_MP913 N$14023 SK2 N$14014 VDD p l=2e-06 w=5e-06
M_MP918 N$14019 N$14015 N$14012 VDD p l=2e-06 w=5e-06
M_MP917 N$14021 SK2 N$14012 VDD p l=2e-06 w=5e-06
M_MP882 0 N$14037 N$14033 VDD p l=2e-06 w=5e-06
M_MP881 0 N$14040 N$14033 VDD p l=2e-06 w=5e-06
M_MP887 P3 N$14040 N$14029 VDD p l=2e-06 w=5e-06
M_MP886 0 N$14037 N$14030 VDD p l=2e-06 w=5e-06
M_MP885 P4 N$14040 N$14030 VDD p l=2e-06 w=5e-06
M_MP229 N$1180 N$14095 N$266 VDD p l=2e-06 w=5e-06
M_MP357 N$372 N$14096 N$386 VDD p l=2e-06 w=5e-06
M_MP379 N$11787 N$11790 VDD VDD p l=2e-06 w=6e-06
M_MP384 N$11779 N$11778 VDD VDD p l=2e-06 w=6e-06
M_MP376 N$11783 N$11789 N$11790 VDD p l=2e-06 w=6e-06
M_MP893 N$14039 SK1 N$14025 VDD p l=2e-06 w=5e-06
M_MP892 0 N$14037 N$14027 VDD p l=2e-06 w=5e-06
M_MP932 N$14013 SK3 N$14004 VDD p l=2e-06 w=5e-06
M_MP937 N$14008 N$14006 N$14002 VDD p l=2e-06 w=5e-06
M_MP936 N$14011 SK3 N$14002 VDD p l=2e-06 w=5e-06
M_MP935 N$14009 N$14006 N$14003 VDD p l=2e-06 w=5e-06
M_MP750 N$11335 N$11332 VDD VDD p l=2e-06 w=6e-06
M_MP10 N$14 N$2 VDD VDD p l=2e-06 w=6e-06
M_MP9 N$13 N$8 VDD VDD p l=2e-06 w=6e-06
M_MP505 N$12429 N$12633 VDD VDD p l=2e-06 w=6e-06
M_MP502 N$1571 N$1570 VDD VDD p l=2e-06 w=6e-06
M_MP517 N$1559 N$1558 VDD VDD p l=2e-06 w=5e-06
M_MP2 N$2 add_one VDD VDD p l=2e-06 w=6e-06
M_MP1 N$2 N$3 VDD VDD p l=2e-06 w=6e-06
M_MP742 N$11331 N$11330 VDD VDD p l=2e-06 w=6e-06
M_MP754 N$382 N$11337 VDD VDD p l=2e-06 w=6e-06
M_MP241 N$279 N$385 VDD VDD p l=2e-06 w=6e-06
M_MP405 N$1180 N$1177 VDD VDD p l=2e-06 w=5e-06
M_MP323 N$310 N$11347 N$14086 VDD p l=2e-06 w=5e-06
M_MP403 N$1176 N$1179 VDD VDD p l=2e-06 w=5e-06
M_MP404 N$1177 0 N$1176 VDD p l=2e-06 w=5e-06
M_MP19 N$25 N$20 VDD VDD p l=2e-06 w=6e-06
M_MP18 N$22 N$17 VDD VDD p l=2e-06 w=6e-06
M_MP17 N$21 N$16 VDD VDD p l=2e-06 w=6e-06
M_MP254 N$301 N$298 VDD VDD p l=2e-06 w=6e-06
M_MP196 N$222 N$207 N$219 VDD p l=2e-06 w=3e-06
M_MP150 N$166 N$162 VDD VDD p l=2e-06 w=3e-06
M_MP368 0 N$409 N$394 VDD p l=2e-06 w=5e-06
M_MP367 N$412 N$14096 N$392 VDD p l=2e-06 w=5e-06
M_MP366 0 N$409 N$392 VDD p l=2e-06 w=5e-06
M_MP447 N$12835 N$1627 VDD VDD p l=2e-06 w=3e-06
M_MP449 N$1622 N$1620 VDD VDD p l=2e-06 w=3e-06
M_MP369 N$397 N$14096 N$394 VDD p l=2e-06 w=5e-06
M_MP448 N$1622 N$1599 VDD VDD p l=2e-06 w=3e-06
M_MP6 N$8 add_one N$7 VDD p l=2e-06 w=6e-06
M_MP96 N$96 N$386 VDD VDD p l=2e-06 w=3e-06
M_MP95 N$96 0 VDD VDD p l=2e-06 w=3e-06
M_MP228 N$1179 N$265 N$266 VDD p l=2e-06 w=5e-06
M_MP98 N$100 N$84 N$96 VDD p l=2e-06 w=3e-06
M_MP305 N$334 CK VDD VDD p l=2e-06 w=5e-06
M_MP518 N$1557 N$11083 N$1559 VDD p l=2e-06 w=5e-06
M_MP267 N$310 N$311 VDD VDD p l=2e-06 w=6e-06
M_MP61 N$271 CK N$282 VDD p l=2e-06 w=6e-06
M_MP269 N$306 CK VDD VDD p l=2e-06 w=5e-06
M_MP268 N$311 N$309 VDD VDD p l=2e-06 w=6e-06
M_MP450 N$1619 N$1620 N$1622 VDD p l=2e-06 w=3e-06
M_MP8 N$10 add_one VDD VDD p l=2e-06 w=6e-06
M_MP333 N$345 N$11347 N$14091 VDD p l=2e-06 w=5e-06
M_MP370 0 N$409 N$395 VDD p l=2e-06 w=5e-06
M_MP334 OUT8 N$11347 N$398 VDD p l=2e-06 w=5e-06
M_MP311 N$344 CK N$345 VDD p l=2e-06 w=6e-06
M_MP310 N$342 N$341 N$344 VDD p l=2e-06 w=6e-06
M_MP252 N$242 CK N$298 VDD p l=2e-06 w=6e-06
M_MP178 N$200 N$196 VDD VDD p l=2e-06 w=3e-06
M_MP107 N$108 N$100 N$105 VDD p l=2e-06 w=3e-06
M_MP135 N$144 N$136 N$141 VDD p l=2e-06 w=3e-06
M_MP134 N$144 N$120 N$143 VDD p l=2e-06 w=3e-06
M_MP133 N$143 N$388 N$142 VDD p l=2e-06 w=3e-06
M_MP132 N$142 0 N$141 VDD p l=2e-06 w=3e-06
M_MP176 N$196 N$173 N$195 VDD p l=2e-06 w=3e-06
M_MP773 N$12429 RST N$1599 VDD p l=2e-06 w=5e-06
M_MP772 0 N$11813 N$1599 VDD p l=2e-06 w=5e-06
M_MP771 N$11794 B0 VDD VDD p l=2e-06 w=3e-06
M_MP354 N$398 N$14096 N$385 VDD p l=2e-06 w=5e-06
M_MP165 N$185 N$14079 VDD VDD p l=2e-06 w=3e-06
M_MP166 N$185 N$392 VDD VDD p l=2e-06 w=3e-06
M_MP314 N$341 CK VDD VDD p l=2e-06 w=5e-06
M_MP149 N$162 N$154 N$159 VDD p l=2e-06 w=3e-06
M_MP148 N$162 N$138 N$161 VDD p l=2e-06 w=3e-06
M_MP147 N$161 N$389 N$160 VDD p l=2e-06 w=3e-06
M_MP205 N$230 N$222 N$227 VDD p l=2e-06 w=3e-06
M_MP155 N$171 N$14078 N$170 VDD p l=2e-06 w=3e-06
M_MP154 N$171 N$156 N$168 VDD p l=2e-06 w=3e-06
M_MP123 N$132 0 VDD VDD p l=2e-06 w=3e-06
M_MP285 N$324 N$325 VDD VDD p l=2e-06 w=6e-06
M_MP284 N$323 CK N$324 VDD p l=2e-06 w=6e-06
M_MP62 N$282 N$283 N$286 VDD p l=2e-06 w=6e-06
M_MP180 N$202 N$394 VDD VDD p l=2e-06 w=3e-06
M_MP179 N$202 N$14080 VDD VDD p l=2e-06 w=3e-06
M_MP689 N$14098 CK VDD VDD p l=2e-06 w=5e-06
M_MP644 N$1437 N$1441 VDD VDD p l=2e-06 w=3e-06
M_MP681 N$14097 CK N$1406 VDD p l=2e-06 w=6e-06
M_MP175 N$195 N$392 N$194 VDD p l=2e-06 w=3e-06
M_MP174 N$194 N$14079 N$193 VDD p l=2e-06 w=3e-06
M_MP173 N$193 N$392 VDD VDD p l=2e-06 w=3e-06
M_MP202 N$228 N$14081 N$227 VDD p l=2e-06 w=3e-06
M_MP65 N$286 N$283 N$288 VDD p l=2e-06 w=6e-06
M_MP286 N$325 N$323 VDD VDD p l=2e-06 w=6e-06
M_MP301 N$335 N$334 N$337 VDD p l=2e-06 w=6e-06
M_MP300 N$335 N$336 VDD VDD p l=2e-06 w=6e-06
M_MP251 N$292 CK VDD VDD p l=2e-06 w=5e-06
M_MP195 N$221 N$395 N$219 VDD p l=2e-06 w=3e-06
M_MP194 N$219 N$395 VDD VDD p l=2e-06 w=3e-06
M_MP193 N$219 N$14081 VDD VDD p l=2e-06 w=3e-06
M_MP255 N$300 N$301 VDD VDD p l=2e-06 w=6e-06
M_MP849 N$13965 N$14005 VDD VDD p l=2e-06 w=3e-06
M_MP848 N$13965 N$14090 VDD VDD p l=2e-06 w=3e-06
M_MP875 OUT7 N$13991 VDD VDD p l=2e-06 w=3e-06
M_MP204 N$230 N$207 N$229 VDD p l=2e-06 w=3e-06
M_MP203 N$229 N$395 N$228 VDD p l=2e-06 w=3e-06
M_MP225 N$217 N$265 N$262 VDD p l=2e-06 w=5e-06
M_MP67 N$361 N$290 VDD VDD p l=2e-06 w=6e-06
M_MP66 N$288 CK N$361 VDD p l=2e-06 w=6e-06
M_MP207 N$112 N$265 N$237 VDD p l=2e-06 w=5e-06
M_MP713 N$1384 CK N$14092 VDD p l=2e-06 w=6e-06
M_MP686 N$1402 CK N$14046 VDD p l=2e-06 w=6e-06
M_MP685 N$1404 N$14098 N$1402 VDD p l=2e-06 w=6e-06
M_MP690 N$1410 CK N$1400 VDD p l=2e-06 w=6e-06
M_MP164 N$183 N$179 VDD VDD p l=2e-06 w=3e-06
M_MP161 N$178 N$390 N$177 VDD p l=2e-06 w=3e-06
M_MP113 N$118 0 N$117 VDD p l=2e-06 w=3e-06
M_MP112 N$118 N$102 N$114 VDD p l=2e-06 w=3e-06
M_MP111 N$117 N$387 N$114 VDD p l=2e-06 w=3e-06
M_MP680 0 N$1557 N$1408 VDD p l=2e-06 w=5e-06
M_MP880 0 N$14037 N$14035 VDD p l=2e-06 w=5e-06
M_MP879 0 N$14040 N$14035 VDD p l=2e-06 w=5e-06
M_MP884 0 N$14037 N$14031 VDD p l=2e-06 w=5e-06
M_MP883 0 N$14040 N$14031 VDD p l=2e-06 w=5e-06
M_MP850 N$13966 N$14005 N$13965 VDD p l=2e-06 w=3e-06
M_MP160 N$177 N$14078 N$176 VDD p l=2e-06 w=3e-06
M_MP159 N$176 N$390 VDD VDD p l=2e-06 w=3e-06
M_MP751 N$11334 N$11335 VDD VDD p l=2e-06 w=6e-06
M_MP735 N$11344 CK N$11326 VDD p l=2e-06 w=6e-06
M_MP734 N$11321 CK VDD VDD p l=2e-06 w=5e-06
M_MP733 N$11325 N$11324 VDD VDD p l=2e-06 w=6e-06
M_MP353 0 N$409 N$385 VDD p l=2e-06 w=5e-06
M_MP359 N$410 N$14096 N$387 VDD p l=2e-06 w=5e-06
M_MP360 P3 N$409 N$388 VDD p l=2e-06 w=5e-06


*.ends mynand3

* Auxiliary circuit for power analysis
Cp Pav 0 100p
Rp Pav 0 100k
Fp 0 Pav Vtstp 0.003125
*Output load capacitance if you have any

*Cload1 out GND 200fF
.MODEL n NMOS LEVEL = 3
+ TOX = 200E-10 NSUB = 1E17 GAMMA = 0.5
+ PHI = 0.7 VTO = 0.8 DELTA = 3.0
+ UO = 650 ETA = 3.0E-6 THETA = 0.1
+ KP = 120E-6 VMAX = 1E5 KAPPA = 0.3
+ RSH = 0 NFS = 1E12 TPG = 1
+ XJ = 500E-9 LD = 100E-9
+ CGDO = 200E-12 CGSO = 200E-12 CGBO = 1E-10
+ CJ = 400E-6 PB = 1 MJ = 0.5
+ CJSW = 300E-12 MJSW = 0.5

.MODEL p PMOS LEVEL = 3
+ TOX = 200E-10 NSUB = 1E17 GAMMA = 0.6
+ PHI = 0.7 VTO = -0.9 DELTA = 0.1
+ UO = 250 ETA = 0 THETA = 0.1
+ KP = 40E-6 VMAX = 5E4 KAPPA = 1
+ RSH = 0 NFS = 1E12 TPG = -1
+ XJ = 500E-9 LD = 100E-9
+ CGDO = 200E-12 CGSO = 200E-12 CGBO = 1E-10
+ CJ = 400E-6 PB = 1 MJ = 0.5
+ CJSW = 300E-12 MJSW = 0.5

*Define power rails
Vddt top 0 5
Vtstp top Vdd 0
Vss GND 0 0

* Define input voltages of A and B

Vck CK 0 PWL(0 5 20N 5 20.1N 0 40N 0 40.1N 5 60N 5 60.1N 0 80N 0 80.1N 5 100N 5 
+ 100.1N 0 120N 0 120.1N 5 140N 5 140.1N 0 160N 0 160.1N 5 180N 5 180.1N 0 200N 0
+ 200.1N 5 220N 5 220.1N 0 240N 0 240.1N 5 260N 5 260.1N 0 280N 0 280.1N 5 300N 5 
+ 300.1N 0 320N 0 320.1N 5 340N 5 340.1N 0 360N 0 360.1N 5 380N 5 380.1N 0 400N 0 
+ 400.1N 5 420N 5 420.1N 0 440N 0 440.1N 5 460N 5 460.1N 0 480N 0 480.1N 5 500N 5)

Va5 A5 0 PWL(0 5 20N 5 20.1N 5 40N 5 40.1N 5 60N 5 60.1N 5 80N 5 80.1N 5 100N 5 
+ 100.1N 5 120N 5 120.1N 5 140N 5 140.1N 5 160N 5 160.1N 5 180N 5 180.1N 5 200N 5
+ 200.1N 0 220N 0 220.1N 0 240N 0 240.1N 0 260N 0 260.1N 0 280N 0 280.1N 0 300N 0 
+ 300.1N 0 320N 0 320.1N 0 340N 0 340.1N 0 360N 0 360.1N 0 380N 0 380.1N 0 400N 0 
+ 400.1N 0 420N 0 420.1N 0 440N 0 440.1N 0 460N 0 460.1N 0 480N 0 480.1N 0 500N 0)

Vp1 P1 0 PWL(0 5 20N 5 20.1N 5 40N 5 40.1N 5 60N 5 60.1N 5 80N 5 80.1N 5 100N 5 
+ 100.1N 5 120N 5 120.1N 5 140N 5 140.1N 5 160N 5 160.1N 5 180N 5 180.1N 5 200N 5
+ 200.1N 5 220N 5 220.1N 5 240N 5 240.1N 5 260N 5 260.1N 5 280N 5 280.1N 5 300N 5 
+ 300.1N 5 320N 5 320.1N 5 340N 5 340.1N 5 360N 5 360.1N 5 380N 5 380.1N 5 400N 5 
+ 400.1N 5 420N 5 420.1N 5 440N 5 440.1N 5 460N 5 460.1N 5 480N 5 480.1N 5 500N 5)

Vp2 P2 0 PWL(0 0 20N 0 20.1N 0 40N 0 40.1N 0 60N 0 60.1N 0 80N 0 80.1N 0 100N 0 
+ 100.1N 0 120N 0 120.1N 0 140N 0 140.1N 0 160N 0 160.1N 0 180N 0 180.1N 0 200N 0
+ 200.1N 0 220N 0 220.1N 0 240N 0 240.1N 0 260N 0 260.1N 0 280N 0 280.1N 0 300N 0 
+ 300.1N 0 320N 0 320.1N 0 340N 0 340.1N 0 360N 0 360.1N 0 380N 0 380.1N 0 400N 0 
+ 400.1N 0 420N 0 420.1N 0 440N 0 440.1N 0 460N 0 460.1N 0 480N 0 480.1N 0 500N 0)

Vp3 P3 0 PWL(0 5 20N 5 20.1N 5 40N 5 40.1N 5 60N 5 60.1N 5 80N 5 80.1N 5 100N 5 
+ 100.1N 5 120N 5 120.1N 5 140N 5 140.1N 5 160N 5 160.1N 5 180N 5 180.1N 5 200N 5
+ 200.1N 5 220N 5 220.1N 5 240N 5 240.1N 5 260N 5 260.1N 5 280N 5 280.1N 5 300N 5 
+ 300.1N 5 320N 5 320.1N 5 340N 5 340.1N 5 360N 5 360.1N 5 380N 5 380.1N 5 400N 5 
+ 400.1N 5 420N 5 420.1N 5 440N 5 440.1N 5 460N 5 460.1N 5 480N 5 480.1N 5 500N 5)

Vp4 P4 0 PWL(0 0 20N 0 20.1N 0 40N 0 40.1N 0 60N 0 60.1N 0 80N 0 80.1N 0 100N 0 
+ 100.1N 0 120N 0 120.1N 0 140N 0 140.1N 0 160N 0 160.1N 0 180N 0 180.1N 0 200N 0
+ 200.1N 0 220N 0 220.1N 0 240N 0 240.1N 0 260N 0 260.1N 0 280N 0 280.1N 0 300N 0 
+ 300.1N 0 320N 0 320.1N 0 340N 0 340.1N 0 360N 0 360.1N 0 380N 0 380.1N 0 400N 0 
+ 400.1N 0 420N 0 420.1N 0 440N 0 440.1N 0 460N 0 460.1N 0 480N 0 480.1N 0 500N 0)

Vrst RST 0 PWL(0 5 20N 5 20.1N 5 40N 5 40.1N 0 60N 0 60.1N 0 80N 0 80.1N 0 100N 0 
+ 100.1N 0 120N 0 120.1N 0 140N 0 140.1N 0 160N 0 160.1N 0 180N 0 180.1N 0 200N 0
+ 200.1N 0 220N 0 220.1N 0 240N 0 240.1N 0 260N 0 260.1N 0 280N 0 280.1N 0 300N 0 
+ 300.1N 0 320N 0 320.1N 0 340N 0 340.1N 0 360N 0 360.1N 0 380N 0 380.1N 0 400N 0 
+ 400.1N 0 420N 0 420.1N 0 440N 0 440.1N 0 460N 0 460.1N 0 480N 0 480.1N 0 500N 0)

Vb0 B0 0 PWL(0 5 20N 5 20.1N 5 40N 5 40.1N 5 60N 5 60.1N 5 80N 5 80.1N 5 100N 5 
+ 100.1N 5 120N 5 120.1N 5 140N 5 140.1N 5 160N 5 160.1N 5 180N 5 180.1N 5 200N 5
+ 200.1N 5 220N 5 220.1N 5 240N 5 240.1N 5 260N 5 260.1N 5 280N 5 280.1N 5 300N 5 
+ 300.1N 5 320N 5 320.1N 5 340N 5 340.1N 5 360N 5 360.1N 5 380N 5 380.1N 5 400N 5 
+ 400.1N 5 420N 5 420.1N 5 440N 5 440.1N 5 460N 5 460.1N 5 480N 5 480.1N 5 500N 5)

Vb1 B1 0 PWL(0 0 20N 0 20.1N 0 40N 0 40.1N 0 60N 0 60.1N 0 80N 0 80.1N 0 100N 0 
+ 100.1N 0 120N 0 120.1N 0 140N 0 140.1N 0 160N 0 160.1N 0 180N 0 180.1N 0 200N 0
+ 200.1N 0 220N 0 220.1N 0 240N 0 240.1N 0 260N 0 260.1N 0 280N 0 280.1N 0 300N 0 
+ 300.1N 0 320N 0 320.1N 0 340N 0 340.1N 0 360N 0 360.1N 0 380N 0 380.1N 0 400N 0 
+ 400.1N 0 420N 0 420.1N 0 440N 0 440.1N 0 460N 0 460.1N 0 480N 0 480.1N 0 500N 0)

Vb2 B2 0 PWL(0 5 20N 5 20.1N 5 40N 5 40.1N 5 60N 5 60.1N 5 80N 5 80.1N 5 100N 5 
+ 100.1N 5 120N 5 120.1N 5 140N 5 140.1N 5 160N 5 160.1N 5 180N 5 180.1N 5 200N 5
+ 200.1N 5 220N 5 220.1N 5 240N 5 240.1N 5 260N 5 260.1N 5 280N 5 280.1N 5 300N 5 
+ 300.1N 5 320N 5 320.1N 5 340N 5 340.1N 5 360N 5 360.1N 5 380N 5 380.1N 5 400N 5 
+ 400.1N 5 420N 5 420.1N 5 440N 5 440.1N 5 460N 5 460.1N 5 480N 5 480.1N 5 500N 5)

Vb3 B3 0 PWL(0 0 20N 0 20.1N 0 40N 0 40.1N 0 60N 0 60.1N 0 80N 0 80.1N 0 100N 0 
+ 100.1N 0 120N 0 120.1N 0 140N 0 140.1N 0 160N 0 160.1N 0 180N 0 180.1N 0 200N 0
+ 200.1N 0 220N 0 220.1N 0 240N 0 240.1N 0 260N 0 260.1N 0 280N 0 280.1N 0 300N 0 
+ 300.1N 0 320N 0 320.1N 0 340N 0 340.1N 0 360N 0 360.1N 0 380N 0 380.1N 0 400N 0 
+ 400.1N 0 420N 0 420.1N 0 440N 0 440.1N 0 460N 0 460.1N 0 480N 0 480.1N 0 500N 0)

Vc C 0 PWL(0 5 20N 5 20.1N 5 40N 5 40.1N 5 60N 5 60.1N 5 80N 5 80.1N 5 100N 5 
+ 100.1N 5 120N 5 120.1N 5 140N 5 140.1N 5 160N 5 160.1N 5 180N 5 180.1N 5 200N 5
+ 200.1N 5 220N 5 220.1N 5 240N 5 240.1N 5 260N 5 260.1N 5 280N 5 280.1N 5 300N 5 
+ 300.1N 5 320N 5 320.1N 5 340N 5 340.1N 5 360N 5 360.1N 5 380N 5 380.1N 5 400N 5 
+ 400.1N 5 420N 5 420.1N 5 440N 5 440.1N 5 460N 5 460.1N 5 480N 5 480.1N 5 500N 5)

Vadd_one add_one 0 PWL(0 5 20N 5 20.1N 5 40N 5 40.1N 5 60N 5 60.1N 5 80N 5 80.1N 5 100N 5 
+ 100.1N 5 120N 5 120.1N 5 140N 5 140.1N 5 160N 5 160.1N 5 180N 5 180.1N 5 200N 5
+ 200.1N 5 220N 5 220.1N 5 240N 5 240.1N 5 260N 5 260.1N 5 280N 5 280.1N 5 300N 5 
+ 300.1N 5 320N 5 320.1N 5 340N 5 340.1N 5 360N 5 360.1N 5 380N 5 380.1N 5 400N 5 
+ 400.1N 5 420N 5 420.1N 5 440N 5 440.1N 5 460N 5 460.1N 5 480N 5 480.1N 5 500N 5)


*Define transient simulation and probe voltage/current signals
.TRAN 20N 500N
.PROBE V(*) I(*)
.end
 



