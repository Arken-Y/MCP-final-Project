




*.subckt mynand3 A B GND Out Vdd



* MAIN CELL: Component pathname : /home/mentor/jack/jaggu
*
        MP142 N$707 N$1055 VDD VDD p L=2u W=6u
        MN142 N$707 N$1055 GND GND n L=2u W=6u
        MP76 N$1034 N$6186 VDD VDD p L=2u W=6u
        MN75 N$1034 N$6186 N$1030 GND n L=2u W=6u
        MP75 N$1034 N$4991 VDD VDD p L=2u W=6u
        MN74 N$37 N$1032 GND GND n L=2u W=6u
        MP74 N$37 N$1032 VDD VDD p L=2u W=6u
        MN276 N$4348 N$4352 GND GND n L=2u W=6u
        MP276 N$4348 N$4352 VDD VDD p L=2u W=6u
        MP275 N$4349 CK N$4348 VDD p L=2u W=6u
        MN275 N$4348 N$4354 N$4349 GND n L=2u W=6u
        MP274 N$4350 N$4354 N$4349 VDD p L=2u W=6u
        MN274 N$4349 CK N$4350 GND n L=2u W=6u
        MN273 N$4350 N$4353 GND GND n L=2u W=6u
        MP273 N$4350 N$4353 VDD VDD p L=2u W=6u
        MN272 N$4353 N$4351 GND GND n L=2u W=6u
        MP272 N$4353 N$4351 VDD VDD p L=2u W=6u
        MP271 N$4351 N$4354 N$4350 VDD p L=2u W=6u
        MN271 N$4350 CK N$4351 GND n L=2u W=6u
        MP270 N$4320 CK N$4351 VDD p L=2u W=6u
        MN113 N$947 N$2908 GND GND n L=2u W=3u
        MN112 N$948 N$2908 GND GND n L=2u W=3u
        MN111 N$945 N$41 N$947 GND n L=2u W=3u
        MN110 N$947 N$1579 GND GND n L=2u W=3u
        MN109 N$946 N$945 GND GND n L=2u W=3u
        MP113 N$945 N$1579 N$944 VDD p L=2u W=3u
        MP112 N$945 N$41 N$943 VDD p L=2u W=3u
        MP111 N$944 N$2908 N$943 VDD p L=2u W=3u
        MP110 N$943 N$2908 VDD VDD p L=2u W=3u
        MP109 N$943 N$1579 VDD VDD p L=2u W=3u
        MN114 N$945 N$1579 N$948 GND n L=2u W=3u
        MP191 N$1014 N$1607 VDD VDD p L=2u W=3u
        MP192 N$1014 N$1584 VDD VDD p L=2u W=3u
        MP533 N$5423 N$5422 VDD VDD p L=2u W=6u
        MN532 N$5422 N$5427 GND GND n L=2u W=6u
        MP532 N$5422 N$5427 VDD VDD p L=2u W=6u
        MP531 N$5427 N$5426 N$5423 VDD p L=2u W=6u
        MN531 N$5423 CK N$5427 GND n L=2u W=6u
        MP530 N$5430 CK N$5427 VDD p L=2u W=6u
        MN530 N$5427 N$5426 N$5430 GND n L=2u W=6u
        MN493 N$5453 N$5458 GND GND n L=2u W=3u
        MN492 N$5456 N$5471 N$5454 GND n L=2u W=3u
        MN491 N$5454 N$5459 GND GND n L=2u W=3u
        MP502 N$5449 N$5456 N$5452 VDD p L=2u W=3u
        MP501 N$5449 N$5471 N$5450 VDD p L=2u W=3u
        MP500 N$5450 N$5458 N$5451 VDD p L=2u W=3u
        MP499 N$5451 N$5459 N$5452 VDD p L=2u W=3u
        MP498 N$5452 N$5458 VDD VDD p L=2u W=3u
        MP497 N$5452 N$5459 VDD VDD p L=2u W=3u
        MP496 N$5452 N$5471 VDD VDD p L=2u W=3u
        MN502 N$5449 N$5471 N$5447 GND n L=2u W=3u
        MN501 N$5449 N$5456 N$5448 GND n L=2u W=3u
        MN500 N$5446 N$5458 GND GND n L=2u W=3u
        MN499 N$5447 N$5459 N$5446 GND n L=2u W=3u
        MN498 N$5448 N$5471 GND GND n L=2u W=3u
        MN497 N$5448 N$5458 GND GND n L=2u W=3u
        MN496 N$5448 N$5459 GND GND n L=2u W=3u
        MP505 N$5491 B2 VDD VDD p L=2u W=3u
        MN504 N$5510 B1 GND GND n L=2u W=3u
        MP504 N$5510 B1 VDD VDD p L=2u W=3u
        MP527 N$5511 N$5455 N$5431 VDD p L=2u W=5u
        MN503 N$5445 N$5449 GND GND n L=2u W=3u
        MP1070 N$5224 N$5223 VDD VDD p L=2u W=6u
        MN1076 N$5225 CK GND GND n L=2u W=5u
        MP1075 N$5225 CK VDD VDD p L=2u W=5u
        MN1075 N$5221 N$5222 GND GND n L=2u W=6u
        MP1074 N$5221 N$5222 VDD VDD p L=2u W=6u
        MN55 N$3670 GND N$3672 GND n L=2u W=3u
        MN54 N$3670 N$3664 N$3671 GND n L=2u W=3u
        MN53 N$3673 N$3701 GND GND n L=2u W=3u
        MP36 N$44 N$2904 VDD VDD p L=2u W=3u
        MP35 N$44 GND VDD VDD p L=2u W=3u
        MP34 N$41 N$40 VDD VDD p L=2u W=3u
        MN38 N$49 N$2904 N$50 GND n L=2u W=3u
        MN37 N$48 GND GND GND n L=2u W=3u
        MN36 N$48 N$2906 GND GND n L=2u W=3u
        MN35 N$48 N$2904 GND GND n L=2u W=3u
        MP41 N$47 N$40 N$44 VDD p L=2u W=3u
        MN447 N$5505 N$5508 GND GND n L=2u W=3u
        MP451 N$5508 N$5511 N$5509 VDD p L=2u W=3u
        MP450 N$5508 N$5507 N$5512 VDD p L=2u W=3u
        MP449 N$5509 N$5510 N$5512 VDD p L=2u W=3u
        MP448 N$5512 N$5510 VDD VDD p L=2u W=3u
        MP136 N$3704 N$3683 VDD VDD p L=2u W=3u
        MN136 N$3704 N$3683 GND GND n L=2u W=3u
        MP149 N$3687 N$1017 VDD VDD p L=2u W=3u
        MP150 N$3687 N$3456 VDD VDD p L=2u W=3u
        MP151 N$3688 N$3456 N$3687 VDD p L=2u W=3u
        MP152 N$3689 N$3460 N$3687 VDD p L=2u W=3u
        MP195 N$1016 N$1607 N$1015 VDD p L=2u W=3u
        MP193 N$1015 N$1584 N$1014 VDD p L=2u W=3u
        MP194 N$1016 N$946 N$1014 VDD p L=2u W=3u
        MP346 N$5909 N$5357 N$5922 VDD p L=2u W=5u
        MN356 N$5926 N$5357 N$5917 GND n L=2u W=5u
        MN345 N$5920 N$5979 GND GND n L=2u W=5u
        MP345 GND N$5958 N$5920 VDD p L=2u W=5u
        MN344 N$5920 N$5958 A0 GND n L=2u W=5u
        MN1090 N$5210 N$5216 N$5209 GND n L=2u W=3u
        MN1089 N$5207 N$5218 GND GND n L=2u W=3u
        MN1088 N$5208 N$5429 N$5207 GND n L=2u W=3u
        MN1091 N$5210 C N$5208 GND n L=2u W=3u
        MP1094 N$5406 RST N$5459 VDD p L=2u W=5u
        MN1094 N$5459 RST GND GND n L=2u W=5u
        MP1093 GND N$5385 N$5459 VDD p L=2u W=5u
        MP1066 N$5232 CK VDD VDD p L=2u W=5u
        MN1066 N$5227 N$5228 GND GND n L=2u W=6u
        MP1065 N$5227 N$5228 VDD VDD p L=2u W=6u
        MN1065 N$5383 N$5227 GND GND n L=2u W=6u
        MP1064 N$5383 N$5227 VDD VDD p L=2u W=6u
        MP1063 N$5228 CK N$5383 VDD p L=2u W=6u
        MN1070 N$5223 N$5226 GND GND n L=2u W=6u
        MP1069 N$5223 N$5226 VDD VDD p L=2u W=6u
        MP1068 N$5226 N$5225 N$5224 VDD p L=2u W=6u
        MN1069 N$5224 CK N$5226 GND n L=2u W=6u
        MP1067 N$5432 CK N$5226 VDD p L=2u W=6u
        MN1068 N$5226 N$5225 N$5432 GND n L=2u W=6u
        MN1067 N$5232 CK GND GND n L=2u W=5u
        MP1072 N$5222 CK N$5381 VDD p L=2u W=6u
        MN1073 N$5381 N$5225 N$5222 GND n L=2u W=6u
        MP1071 N$5224 N$5225 N$5222 VDD p L=2u W=6u
        MN1072 N$5222 CK N$5224 GND n L=2u W=6u
        MN1071 N$5224 N$5223 GND GND n L=2u W=6u
        MN335 N$5914 N$5979 GND GND n L=2u W=5u
        MP335 GND N$5958 N$5914 VDD p L=2u W=5u
        MN334 N$5914 N$5958 GND GND n L=2u W=5u
        MP334 GND N$5979 N$5914 VDD p L=2u W=5u
        MN433 N$5948 N$5941 N$5939 GND n L=2u W=5u
        MP434 GND N$5941 N$5948 VDD p L=2u W=5u
        MN333 N$5912 N$5979 GND GND n L=2u W=5u
        MN302 N$4315 N$4372 N$4367 GND n L=2u W=6u
        MP301 N$4368 N$4372 N$4367 VDD p L=2u W=6u
        MN451 N$5504 N$5510 GND GND n L=2u W=3u
        MN450 N$5503 N$5510 GND GND n L=2u W=3u
        MN449 N$5508 N$5507 N$5504 GND n L=2u W=3u
        MN448 N$5504 N$5511 GND GND n L=2u W=3u
        MN280 N$4356 CK N$4357 GND n L=2u W=6u
        MP302 N$4367 CK N$4315 VDD p L=2u W=6u
        MP356 N$5917 N$5923 N$5926 VDD p L=2u W=5u
        MN355 N$5926 N$5923 N$5916 GND n L=2u W=5u
        MP355 N$5916 N$5357 N$5926 VDD p L=2u W=5u
        MN354 N$5925 N$5357 N$5916 GND n L=2u W=5u
        MP354 N$5916 N$5923 N$5925 VDD p L=2u W=5u
        MN353 N$5925 N$5923 N$5914 GND n L=2u W=5u
        MP353 N$5914 N$5357 N$5925 VDD p L=2u W=5u
        MN350 N$5924 N$5357 N$5914 GND n L=2u W=5u
        MP350 N$5914 N$5923 N$5924 VDD p L=2u W=5u
        MN349 N$5924 N$5923 N$5912 GND n L=2u W=5u
        MP349 N$5912 N$5357 N$5924 VDD p L=2u W=5u
        MN348 N$5923 N$5357 GND GND n L=2u W=5u
        MP348 N$5923 N$5357 VDD VDD p L=2u W=5u
        MN347 N$5922 N$5357 N$5912 GND n L=2u W=5u
        MP347 N$5912 N$5923 N$5922 VDD p L=2u W=5u
        MN346 N$5922 N$5923 N$5909 GND n L=2u W=5u
        MP390 N$5775 GND N$5774 VDD p L=2u W=3u
        MP389 N$5774 N$5948 N$5773 VDD p L=2u W=3u
        MP388 N$5773 N$4322 N$5772 VDD p L=2u W=3u
        MP387 N$5772 N$5948 VDD VDD p L=2u W=3u
        MP386 N$5772 N$4322 VDD VDD p L=2u W=3u
        MP385 N$5772 GND VDD VDD p L=2u W=3u
        MN389 N$5778 N$5948 GND GND n L=2u W=3u
        MN388 N$5777 N$4322 N$5778 GND n L=2u W=3u
        MN387 N$5776 GND GND GND n L=2u W=3u
        MN386 N$5776 N$5948 GND GND n L=2u W=3u
        MN432 N$5951 N$5341 GND GND n L=2u W=5u
        MP432 GND N$5941 N$5951 VDD p L=2u W=5u
        MN431 N$5951 N$5941 N$5938 GND n L=2u W=5u
        MP431 N$5938 N$5341 N$5951 VDD p L=2u W=5u
        MN430 N$5945 N$5341 GND GND n L=2u W=5u
        MP430 GND N$5941 N$5945 VDD p L=2u W=5u
        MN429 N$5945 N$5941 N$5937 GND n L=2u W=5u
        MP429 N$5937 N$5341 N$5945 VDD p L=2u W=5u
        MN428 N$5955 N$5341 N$5939 GND n L=2u W=5u
        MP428 N$5939 N$5941 N$5955 VDD p L=2u W=5u
        MN427 N$5955 N$5941 N$5936 GND n L=2u W=5u
        MP427 N$5936 N$5341 N$5955 VDD p L=2u W=5u
        MN426 N$5896 N$5341 N$5938 GND n L=2u W=5u
        MP426 N$5938 N$5941 N$5896 VDD p L=2u W=5u
        MN425 N$5896 N$5941 N$5935 GND n L=2u W=5u
        MP425 N$5935 N$5341 N$5896 VDD p L=2u W=5u
        MP379 N$5764 N$4322 VDD VDD p L=2u W=3u
        MP433 N$5939 N$5341 N$5948 VDD p L=2u W=5u
        MN337 N$5916 N$5979 GND GND n L=2u W=5u
        MP337 GND N$5958 N$5916 VDD p L=2u W=5u
        MN336 N$5916 N$5958 GND GND n L=2u W=5u
        MP336 GND N$5979 N$5916 VDD p L=2u W=5u
        MP187 N$1008 N$956 N$1007 VDD p L=2u W=3u
        MN66 N$1049 N$6187 N$1050 GND n L=2u W=6u
        MP62 N$4109 N$1043 VDD VDD p L=2u W=6u
        MP68 N$2908 N$1049 VDD VDD p L=2u W=6u
        MN305 N$4372 CK GND GND n L=2u W=5u
        MP305 N$4372 CK VDD VDD p L=2u W=5u
        MN304 N$4370 N$4367 GND GND n L=2u W=6u
        MP304 N$4370 N$4367 VDD VDD p L=2u W=6u
        MN303 N$4315 N$4370 GND GND n L=2u W=6u
        MP303 N$4315 N$4370 VDD VDD p L=2u W=6u
        MN332 N$5912 N$5958 GND GND n L=2u W=5u
        MP332 GND N$5979 N$5912 VDD p L=2u W=5u
        MN331 N$5958 N$5979 GND GND n L=2u W=5u
        MP331 N$5958 N$5979 VDD VDD p L=2u W=5u
        MP333 GND N$5958 N$5912 VDD p L=2u W=5u
        MN330 N$5909 N$5979 GND GND n L=2u W=5u
        MP330 GND N$5958 N$5909 VDD p L=2u W=5u
        MN329 N$5909 N$5958 GND GND n L=2u W=5u
        MP329 GND N$5979 N$5909 VDD p L=2u W=5u
        MP340 A2 N$5979 N$5918 VDD p L=2u W=5u
        MN339 N$5917 N$5979 GND GND n L=2u W=5u
        MP339 GND N$5958 N$5917 VDD p L=2u W=5u
        MN338 N$5917 N$5958 A3 GND n L=2u W=5u
        MP338 A3 N$5979 N$5917 VDD p L=2u W=5u
        MP384 N$5769 N$5766 VDD VDD p L=2u W=3u
        MN384 N$5766 N$4322 N$5771 GND n L=2u W=3u
        MN383 N$5770 N$5948 GND GND n L=2u W=3u
        MN382 N$5771 N$5948 GND GND n L=2u W=3u
        MN381 N$5766 GND N$5770 GND n L=2u W=3u
        MN380 N$5770 N$4322 GND GND n L=2u W=3u
        MN379 N$5769 N$5766 GND GND n L=2u W=3u
        MP1102 GND N$5910 N$5204 VDD p L=2u W=5u
        MN1102 N$5204 N$5910 A2 GND n L=2u W=5u
        MP1101 A2 N$5201 N$5204 VDD p L=2u W=5u
        MN1101 N$6187 N$5201 GND GND n L=2u W=5u
        MP1100 GND N$5910 N$6187 VDD p L=2u W=5u
        MN1105 N$5744 N$5201 GND GND n L=2u W=5u
        MP1104 GND N$5910 N$5744 VDD p L=2u W=5u
        MN1104 N$5744 N$5910 A3 GND n L=2u W=5u
        MP1103 A3 N$5201 N$5744 VDD p L=2u W=5u
        MP1096 A0 N$5201 N$6186 VDD p L=2u W=5u
        MN183 N$1010 N$2902 GND GND n L=2u W=3u
        MP189 N$1009 N$1002 N$1006 VDD p L=2u W=3u
        MP82 N$914 N$1601 VDD VDD p L=2u W=3u
        MP81 N$914 N$707 VDD VDD p L=2u W=3u
        MN89 N$925 N$9 GND GND n L=2u W=3u
        MN108 N$942 N$938 GND GND n L=2u W=3u
        MP108 N$942 N$938 VDD VDD p L=2u W=3u
        MP226 N$5965 N$5966 N$5967 VDD p L=2u W=6u
        MN226 N$5967 CK N$5965 GND n L=2u W=6u
        MP225 N$5400 CK N$5965 VDD p L=2u W=6u
        MN225 N$5965 N$5966 N$5400 GND n L=2u W=6u
        MP188 N$1009 N$2494 N$1008 VDD p L=2u W=3u
        MN62 N$4109 N$1043 GND GND n L=2u W=6u
        MP453 N$5502 N$5507 VDD VDD p L=2u W=3u
        MP452 N$5505 N$5508 VDD VDD p L=2u W=3u
        MN452 N$5508 N$5511 N$5503 GND n L=2u W=3u
        MP67 N$1049 N$6187 VDD VDD p L=2u W=6u
        MN67 N$1050 N$4989 GND GND n L=2u W=6u
        MN1080 N$5215 N$5429 GND GND n L=2u W=3u
        MN1079 N$5507 N$5216 GND GND n L=2u W=3u
        MP1082 N$5216 N$5429 N$5217 VDD p L=2u W=3u
        MP1081 N$5216 C N$5219 VDD p L=2u W=3u
        MP1080 N$5217 N$5218 N$5219 VDD p L=2u W=3u
        MP1086 N$5213 N$5218 VDD VDD p L=2u W=3u
        MP1085 N$5213 N$5429 VDD VDD p L=2u W=3u
        MP1084 N$5213 C VDD VDD p L=2u W=3u
        MP1083 N$5507 N$5216 VDD VDD p L=2u W=3u
        MN1084 N$5216 N$5429 N$5214 GND n L=2u W=3u
        MN1083 N$5215 N$5218 GND GND n L=2u W=3u
        MN1087 N$5209 C GND GND n L=2u W=3u
        MN1086 N$5209 N$5218 GND GND n L=2u W=3u
        MN1085 N$5209 N$5429 GND GND n L=2u W=3u
        MP1090 N$5210 N$5216 N$5213 VDD p L=2u W=3u
        MP1089 N$5210 C N$5211 VDD p L=2u W=3u
        MP1088 N$5211 N$5218 N$5212 VDD p L=2u W=3u
        MP1087 N$5212 N$5429 N$5213 VDD p L=2u W=3u
        MP1091 N$5441 N$5210 VDD VDD p L=2u W=3u
        MN1093 N$5218 B0 GND GND n L=2u W=3u
        MP1092 N$5218 B0 VDD VDD p L=2u W=3u
        MN1092 N$5441 N$5210 GND GND n L=2u W=3u
        MN1100 N$6187 N$5910 A1 GND n L=2u W=5u
        MP1099 A1 N$5201 N$6187 VDD p L=2u W=5u
        MN1099 N$5201 N$5910 GND GND n L=2u W=5u
        MP1098 N$5201 N$5910 VDD VDD p L=2u W=5u
        MN1098 N$6186 N$5201 GND GND n L=2u W=5u
        MP1097 GND N$5910 N$6186 VDD p L=2u W=5u
        MN1103 N$5204 N$5201 GND GND n L=2u W=5u
        MN998 N$5244 CK GND GND n L=2u W=5u
        MP997 N$5244 CK VDD VDD p L=2u W=5u
        MN997 N$5240 N$5241 GND GND n L=2u W=6u
        MP1002 N$5237 N$5238 N$5235 VDD p L=2u W=6u
        MN1003 N$5235 CK N$5237 GND n L=2u W=6u
        MN1002 N$5237 N$5236 GND GND n L=2u W=6u
        MP1001 N$5237 N$5236 VDD VDD p L=2u W=6u
        MN1001 N$5236 N$5239 GND GND n L=2u W=6u
        MP1000 N$5236 N$5239 VDD VDD p L=2u W=6u
        MP1006 N$5238 CK VDD VDD p L=2u W=5u
        MN1006 N$5234 N$5235 GND GND n L=2u W=6u
        MP1005 N$5234 N$5235 VDD VDD p L=2u W=6u
        MN1005 N$4989 N$5234 GND GND n L=2u W=6u
        MP1004 N$4989 N$5234 VDD VDD p L=2u W=6u
        MP1003 N$5235 CK N$4989 VDD p L=2u W=6u
        MN1004 N$4989 N$5238 N$5235 GND n L=2u W=6u
        MP1060 N$5229 N$5233 VDD VDD p L=2u W=6u
        MP1059 N$5233 N$5232 N$5230 VDD p L=2u W=6u
        MN1060 N$5230 CK N$5233 GND n L=2u W=6u
        MP1058 N$5231 CK N$5233 VDD p L=2u W=6u
        MN1059 N$5233 N$5232 N$5231 GND n L=2u W=6u
        MN1097 N$6186 N$5910 A0 GND n L=2u W=5u
        MP1095 N$5440 N$5445 VDD VDD p L=2u W=5u
        MN1096 N$5437 N$5445 GND GND n L=2u W=5u
        MN1095 N$5459 N$5385 N$5406 GND n L=2u W=5u
        MP1076 N$5429 N$5435 N$5231 VDD p L=2u W=5u
        MN1082 N$5214 N$5218 GND GND n L=2u W=3u
        MN1081 N$5216 C N$5215 GND n L=2u W=3u
        MP981 N$5251 N$5250 N$5249 VDD p L=2u W=6u
        MN982 N$5249 CK N$5251 GND n L=2u W=6u
        MP987 N$5246 N$5247 VDD VDD p L=2u W=6u
        MN987 N$4988 N$5246 GND GND n L=2u W=6u
        MP986 N$4988 N$5246 VDD VDD p L=2u W=6u
        MP985 N$5247 CK N$4988 VDD p L=2u W=6u
        MN986 N$4988 N$5250 N$5247 GND n L=2u W=6u
        MP984 N$5249 N$5250 N$5247 VDD p L=2u W=6u
        MN985 N$5247 CK N$5249 GND n L=2u W=6u
        MN991 N$5243 CK N$5245 GND n L=2u W=6u
        MP989 N$5260 CK N$5245 VDD p L=2u W=6u
        MN990 N$5245 N$5244 N$5260 GND n L=2u W=6u
        MN989 N$5250 CK GND GND n L=2u W=5u
        MP988 N$5250 CK VDD VDD p L=2u W=5u
        MN988 N$5246 N$5247 GND GND n L=2u W=6u
        MN994 N$5241 CK N$5243 GND n L=2u W=6u
        MN993 N$5243 N$5242 GND GND n L=2u W=6u
        MP992 N$5243 N$5242 VDD VDD p L=2u W=6u
        MN992 N$5242 N$5245 GND GND n L=2u W=6u
        MP991 N$5242 N$5245 VDD VDD p L=2u W=6u
        MN1074 N$5381 N$5221 GND GND n L=2u W=6u
        MP1073 N$5381 N$5221 VDD VDD p L=2u W=6u
        MP1079 N$5219 N$5218 VDD VDD p L=2u W=3u
        MP1078 N$5219 N$5429 VDD VDD p L=2u W=3u
        MN1078 N$5231 N$5435 IN7 GND n L=2u W=5u
        MP1077 IN7 N$5455 N$5231 VDD p L=2u W=5u
        MN1077 N$5231 N$5455 N$5429 GND n L=2u W=5u
        MN1000 N$5237 CK N$5239 GND n L=2u W=6u
        MP998 N$5259 CK N$5239 VDD p L=2u W=6u
        MN999 N$5239 N$5238 N$5259 GND n L=2u W=6u
        MN966 N$5261 N$5910 N$5299 GND n L=2u W=5u
        MP965 N$5299 N$5264 N$5261 VDD p L=2u W=5u
        MN971 N$5259 N$5264 GND GND n L=2u W=5u
        MP970 GND N$5910 N$5259 VDD p L=2u W=5u
        MN970 N$5259 N$5910 N$5269 GND n L=2u W=5u
        MP969 N$5269 N$5264 N$5259 VDD p L=2u W=5u
        MN969 N$5260 N$5264 GND GND n L=2u W=5u
        MP974 N$5255 N$5254 VDD VDD p L=2u W=6u
        MN974 N$5254 N$5257 GND GND n L=2u W=6u
        MP973 N$5254 N$5257 VDD VDD p L=2u W=6u
        MP972 N$5257 N$6593 N$5255 VDD p L=2u W=6u
        MN973 N$5255 CK N$5257 GND n L=2u W=6u
        MP971 N$6391 CK N$5257 VDD p L=2u W=6u
        MN972 N$5257 N$6593 N$6391 GND n L=2u W=6u
        MN978 N$4990 N$5252 GND GND n L=2u W=6u
        MP977 N$4990 N$5252 VDD VDD p L=2u W=6u
        MP976 N$5253 CK N$4990 VDD p L=2u W=6u
        MN977 N$4990 N$6593 N$5253 GND n L=2u W=6u
        MP975 N$5255 N$6593 N$5253 VDD p L=2u W=6u
        MN976 N$5253 CK N$5255 GND n L=2u W=6u
        MN1007 N$5238 CK GND GND n L=2u W=5u
        MN1064 N$5383 N$5232 N$5228 GND n L=2u W=6u
        MP1062 N$5230 N$5232 N$5228 VDD p L=2u W=6u
        MN1063 N$5228 CK N$5230 GND n L=2u W=6u
        MN1062 N$5230 N$5229 GND GND n L=2u W=6u
        MP1061 N$5230 N$5229 VDD VDD p L=2u W=6u
        MN1061 N$5229 N$5233 GND GND n L=2u W=6u
        MP983 N$5249 N$5248 VDD VDD p L=2u W=6u
        MN983 N$5248 N$5251 GND GND n L=2u W=6u
        MP982 N$5248 N$5251 VDD VDD p L=2u W=6u
        MN714 N$5267 N$5910 GND GND n L=2u W=5u
        MP715 N$5267 N$5910 VDD VDD p L=2u W=5u
        MN713 N$5370 N$5267 N$5378 GND n L=2u W=5u
        MP714 N$5378 N$5910 N$5370 VDD p L=2u W=5u
        MN712 N$5370 N$5910 N$5337 GND n L=2u W=5u
        MP713 N$5337 N$5267 N$5370 VDD p L=2u W=5u
        MN768 N$5353 N$5910 N$5334 GND n L=2u W=5u
        MP769 N$5334 N$5267 N$5353 VDD p L=2u W=5u
        MN716 N$5361 N$5267 N$5376 GND n L=2u W=5u
        MP768 N$5376 N$5910 N$5361 VDD p L=2u W=5u
        MN715 N$5361 N$5910 N$5335 GND n L=2u W=5u
        MP716 N$5335 N$5267 N$5361 VDD p L=2u W=5u
        MN771 N$5345 N$5267 N$5374 GND n L=2u W=5u
        MP772 N$5374 N$5910 N$5345 VDD p L=2u W=5u
        MN770 N$5345 N$5910 N$5333 GND n L=2u W=5u
        MP771 N$5333 N$5267 N$5345 VDD p L=2u W=5u
        MN769 N$5353 N$5267 N$5375 GND n L=2u W=5u
        MP770 N$5375 N$5910 N$5353 VDD p L=2u W=5u
        MN965 N$5264 N$5910 GND GND n L=2u W=5u
        MP990 N$5245 N$5244 N$5243 VDD p L=2u W=6u
        MP996 N$5240 N$5241 VDD VDD p L=2u W=6u
        MN996 N$4991 N$5240 GND GND n L=2u W=6u
        MP995 N$4991 N$5240 VDD VDD p L=2u W=6u
        MP994 N$5241 CK N$4991 VDD p L=2u W=6u
        MN995 N$4991 N$5244 N$5241 GND n L=2u W=6u
        MP993 N$5243 N$5244 N$5241 VDD p L=2u W=6u
        MP999 N$5239 N$5238 N$5237 VDD p L=2u W=6u
        MP967 N$5284 N$5264 N$5260 VDD p L=2u W=5u
        MN967 N$5261 N$5264 GND GND n L=2u W=5u
        MP966 GND N$5910 N$5261 VDD p L=2u W=5u
        MN698 N$5278 N$5282 GND GND n L=2u W=3u
        MN697 N$5277 N$5282 GND GND n L=2u W=3u
        MN696 N$5280 N$5294 N$5278 GND n L=2u W=3u
        MN695 N$5278 B3 GND GND n L=2u W=3u
        MN694 COUTHK-SK N$5280 GND GND n L=2u W=3u
        MP706 N$5273 N$5294 N$5274 VDD p L=2u W=3u
        MP705 N$5274 N$5282 N$5275 VDD p L=2u W=3u
        MP704 N$5275 B3 N$5276 VDD p L=2u W=3u
        MP703 N$5276 N$5282 VDD VDD p L=2u W=3u
        MP702 N$5276 B3 VDD VDD p L=2u W=3u
        MP701 N$5276 N$5294 VDD VDD p L=2u W=3u
        MN704 N$5270 N$5282 GND GND n L=2u W=3u
        MN703 N$5271 B3 N$5270 GND n L=2u W=3u
        MN702 N$5272 N$5294 GND GND n L=2u W=3u
        MN701 N$5272 N$5282 GND GND n L=2u W=3u
        MN700 N$5272 B3 GND GND n L=2u W=3u
        MP707 N$5273 N$5280 N$5276 VDD p L=2u W=3u
        MN708 N$5329 N$5337 GND GND n L=2u W=3u
        MP709 N$5329 N$5337 VDD VDD p L=2u W=3u
        MN707 N$5269 N$5273 GND GND n L=2u W=3u
        MN975 N$5255 N$5254 GND GND n L=2u W=6u
        MP980 N$5261 CK N$5251 VDD p L=2u W=6u
        MN981 N$5251 N$5250 N$5261 GND n L=2u W=6u
        MN980 N$6593 CK GND GND n L=2u W=5u
        MP979 N$6593 CK VDD VDD p L=2u W=5u
        MN979 N$5252 N$5253 GND GND n L=2u W=6u
        MP978 N$5252 N$5253 VDD VDD p L=2u W=6u
        MN984 N$5249 N$5248 GND GND n L=2u W=6u
        MP711 N$5282 N$5333 VDD VDD p L=2u W=3u
        MN709 N$5312 N$5335 GND GND n L=2u W=3u
        MP710 N$5312 N$5335 VDD VDD p L=2u W=3u
        MN671 N$5294 N$5295 GND GND n L=2u W=3u
        MP685 N$5295 B2 N$5296 VDD p L=2u W=3u
        MP684 N$5295 N$5309 N$5298 VDD p L=2u W=3u
        MP683 N$5296 N$5297 N$5298 VDD p L=2u W=3u
        MP682 N$5298 N$5297 VDD VDD p L=2u W=3u
        MP688 N$5291 B2 VDD VDD p L=2u W=3u
        MP687 N$5291 N$5309 VDD VDD p L=2u W=3u
        MP686 N$5294 N$5295 VDD VDD p L=2u W=3u
        MN685 N$5295 B2 N$5292 GND n L=2u W=3u
        MN684 N$5293 N$5297 GND GND n L=2u W=3u
        MN683 N$5292 N$5297 GND GND n L=2u W=3u
        MN686 N$5287 B2 GND GND n L=2u W=3u
        MP693 N$5288 N$5295 N$5291 VDD p L=2u W=3u
        MP692 N$5288 N$5309 N$5289 VDD p L=2u W=3u
        MP691 N$5289 N$5297 N$5290 VDD p L=2u W=3u
        MP690 N$5290 B2 N$5291 VDD p L=2u W=3u
        MP689 N$5291 N$5297 VDD VDD p L=2u W=3u
        MP694 N$5284 N$5288 VDD VDD p L=2u W=3u
        MN692 N$5288 N$5309 N$5286 GND n L=2u W=3u
        MN691 N$5288 N$5295 N$5287 GND n L=2u W=3u
        MN690 N$5285 N$5297 GND GND n L=2u W=3u
        MP964 N$5264 N$5910 VDD VDD p L=2u W=5u
        MN773 N$6391 N$5264 GND GND n L=2u W=5u
        MP963 GND N$5910 N$6391 VDD p L=2u W=5u
        MN772 N$6391 N$5910 N$5314 GND n L=2u W=5u
        MP773 N$5314 N$5264 N$6391 VDD p L=2u W=5u
        MP968 GND N$5910 N$5260 VDD p L=2u W=5u
        MN968 N$5260 N$5910 N$5284 GND n L=2u W=5u
        MN693 N$5284 N$5288 GND GND n L=2u W=3u
        MP700 COUTHK-SK N$5280 VDD VDD p L=2u W=3u
        MN699 N$5280 B3 N$5277 GND n L=2u W=3u
        MP659 N$5313 N$5312 VDD VDD p L=2u W=3u
        MP658 N$5313 B1 VDD VDD p L=2u W=3u
        MN656 N$5314 N$5318 GND GND n L=2u W=3u
        MP657 N$5314 N$5318 VDD VDD p L=2u W=3u
        MN661 N$5308 N$5312 GND GND n L=2u W=3u
        MN660 N$5307 N$5312 GND GND n L=2u W=3u
        MN659 N$5310 N$5324 N$5308 GND n L=2u W=3u
        MN658 N$5308 B1 GND GND n L=2u W=3u
        MN657 N$5309 N$5310 GND GND n L=2u W=3u
        MP662 N$5310 B1 N$5311 VDD p L=2u W=3u
        MP668 N$5304 N$5312 N$5305 VDD p L=2u W=3u
        MP667 N$5305 B1 N$5306 VDD p L=2u W=3u
        MP666 N$5306 N$5312 VDD VDD p L=2u W=3u
        MP665 N$5306 B1 VDD VDD p L=2u W=3u
        MP664 N$5306 N$5324 VDD VDD p L=2u W=3u
        MP663 N$5309 N$5310 VDD VDD p L=2u W=3u
        MN662 N$5310 B1 N$5307 GND n L=2u W=3u
        MN666 N$5301 B1 N$5300 GND n L=2u W=3u
        MN665 N$5302 N$5324 GND GND n L=2u W=3u
        MN664 N$5302 N$5312 GND GND n L=2u W=3u
        MN663 N$5302 B1 GND GND n L=2u W=3u
        MP708 N$5269 N$5273 VDD VDD p L=2u W=3u
        MN706 N$5273 N$5294 N$5271 GND n L=2u W=3u
        MN705 N$5273 N$5280 N$5272 GND n L=2u W=3u
        MN711 N$5297 N$5334 GND GND n L=2u W=3u
        MP712 N$5297 N$5334 VDD VDD p L=2u W=3u
        MN710 N$5282 N$5333 GND GND n L=2u W=3u
        MN667 N$5300 N$5312 GND GND n L=2u W=3u
        MN682 N$5295 N$5309 N$5293 GND n L=2u W=3u
        MN681 N$5293 B2 GND GND n L=2u W=3u
        MN641 N$5333 N$5910 N$5406 GND n L=2u W=5u
        MP641 N$5406 N$5338 N$5333 VDD p L=2u W=5u
        MN640 N$5334 N$5338 GND GND n L=2u W=5u
        MP640 GND N$5910 N$5334 VDD p L=2u W=5u
        MN643 N$5324 N$5327 GND GND n L=2u W=3u
        MP647 N$5327 B0 N$5328 VDD p L=2u W=3u
        MP646 N$5327 C N$5331 VDD p L=2u W=3u
        MP645 N$5328 N$5329 N$5331 VDD p L=2u W=3u
        MP644 N$5331 N$5329 VDD VDD p L=2u W=3u
        MP643 N$5331 B0 VDD VDD p L=2u W=3u
        MP649 N$5321 C VDD VDD p L=2u W=3u
        MP648 N$5324 N$5327 VDD VDD p L=2u W=3u
        MN648 N$5327 B0 N$5322 GND n L=2u W=3u
        MN647 N$5323 N$5329 GND GND n L=2u W=3u
        MN646 N$5322 N$5329 GND GND n L=2u W=3u
        MN645 N$5327 C N$5323 GND n L=2u W=3u
        MN644 N$5323 B0 GND GND n L=2u W=3u
        MP656 N$5318 N$5327 N$5321 VDD p L=2u W=3u
        MP655 N$5318 C N$5319 VDD p L=2u W=3u
        MP654 N$5319 N$5329 N$5320 VDD p L=2u W=3u
        MP653 N$5320 B0 N$5321 VDD p L=2u W=3u
        MN689 N$5286 B2 N$5285 GND n L=2u W=3u
        MN688 N$5287 N$5309 GND GND n L=2u W=3u
        MN687 N$5287 N$5297 GND GND n L=2u W=3u
        MP699 N$5280 B3 N$5281 VDD p L=2u W=3u
        MP698 N$5280 N$5294 N$5283 VDD p L=2u W=3u
        MP697 N$5281 N$5282 N$5283 VDD p L=2u W=3u
        MP696 N$5283 N$5282 VDD VDD p L=2u W=3u
        MP695 N$5283 B3 VDD VDD p L=2u W=3u
        MN649 N$5317 B0 GND GND n L=2u W=3u
        MP661 N$5310 N$5324 N$5313 VDD p L=2u W=3u
        MP660 N$5311 N$5312 N$5313 VDD p L=2u W=3u
        MP598 N$5370 CK N$5372 VDD p L=2u W=6u
        MN598 N$5372 N$5371 N$5370 GND n L=2u W=6u
        MN597 N$5374 N$5379 GND GND n L=2u W=5u
        MP597 GND N$5387 N$5374 VDD p L=2u W=5u
        MN596 N$5374 N$5387 N$5381 GND n L=2u W=5u
        MP602 N$5368 N$5371 N$5366 VDD p L=2u W=6u
        MN602 N$5366 CK N$5368 GND n L=2u W=6u
        MN601 N$5368 N$5367 GND GND n L=2u W=6u
        MP601 N$5368 N$5367 VDD VDD p L=2u W=6u
        MN600 N$5367 N$5372 GND GND n L=2u W=6u
        MP600 N$5367 N$5372 VDD VDD p L=2u W=6u
        MP599 N$5372 N$5371 N$5368 VDD p L=2u W=6u
        MN605 N$5364 N$5366 GND GND n L=2u W=6u
        MP605 N$5364 N$5366 VDD VDD p L=2u W=6u
        MN604 SK0 N$5364 GND GND n L=2u W=6u
        MP604 SK0 N$5364 VDD VDD p L=2u W=6u
        MP603 N$5366 CK SK0 VDD p L=2u W=6u
        MN603 SK0 N$5371 N$5366 GND n L=2u W=6u
        MP608 N$5363 N$5362 N$5360 VDD p L=2u W=6u
        MN608 N$5360 CK N$5363 GND n L=2u W=6u
        MP651 N$5321 N$5329 VDD VDD p L=2u W=3u
        MP650 N$5321 B0 VDD VDD p L=2u W=3u
        MN655 N$5318 C N$5316 GND n L=2u W=3u
        MN654 N$5318 N$5327 N$5317 GND n L=2u W=3u
        MN653 N$5315 N$5329 GND GND n L=2u W=3u
        MN652 N$5316 B0 N$5315 GND n L=2u W=3u
        MN651 N$5317 C GND GND n L=2u W=3u
        MN650 N$5317 N$5329 GND GND n L=2u W=3u
        MP610 N$5360 N$5359 VDD VDD p L=2u W=6u
        MN609 N$5359 N$5363 GND GND n L=2u W=6u
        MP609 N$5359 N$5363 VDD VDD p L=2u W=6u
        MP582 N$5385 RST VDD VDD p L=2u W=5u
        MN581 N$5429 N$5385 N$5383 GND n L=2u W=5u
        MP581 N$5383 RST N$5429 VDD p L=2u W=5u
        MN580 N$5429 RST A5 GND n L=2u W=5u
        MN586 N$5492 N$5385 N$5413 GND n L=2u W=5u
        MP586 N$5413 RST N$5492 VDD p L=2u W=5u
        MN585 N$5492 RST GND GND n L=2u W=5u
        MP585 GND N$5385 N$5492 VDD p L=2u W=5u
        MN584 N$5511 N$5385 N$5420 GND n L=2u W=5u
        MP584 N$5420 RST N$5511 VDD p L=2u W=5u
        MP590 GND N$5387 N$5378 VDD p L=2u W=5u
        MN589 N$5378 N$5387 N$5383 GND n L=2u W=5u
        MP589 N$5383 N$5379 N$5378 VDD p L=2u W=5u
        MN588 N$5475 N$5385 N$5381 GND n L=2u W=5u
        MP588 N$5381 RST N$5475 VDD p L=2u W=5u
        MN587 N$5475 RST GND GND n L=2u W=5u
        MP587 GND N$5385 N$5475 VDD p L=2u W=5u
        MP593 GND N$5387 N$5376 VDD p L=2u W=5u
        MN592 N$5376 N$5387 N$5420 GND n L=2u W=5u
        MP592 N$5420 N$5379 N$5376 VDD p L=2u W=5u
        MP624 N$5354 CK VDD VDD p L=2u W=5u
        MN623 N$5348 N$5350 GND GND n L=2u W=6u
        MP623 N$5348 N$5350 VDD VDD p L=2u W=6u
        MN622 N$5349 N$5348 GND GND n L=2u W=6u
        MP622 N$5349 N$5348 VDD VDD p L=2u W=6u
        MP621 N$5350 CK N$5349 VDD p L=2u W=6u
        MP627 N$5343 N$5347 VDD VDD p L=2u W=6u
        MP626 N$5347 N$5346 N$5344 VDD p L=2u W=6u
        MP594 N$5413 N$5379 N$5375 VDD p L=2u W=5u
        MN593 N$5376 N$5379 GND GND n L=2u W=5u
        MN599 N$5368 CK N$5372 GND n L=2u W=6u
        MP566 N$5394 CK N$5403 VDD p L=2u W=6u
        MN566 N$5403 N$5397 N$5394 GND n L=2u W=6u
        MP565 N$5396 N$5397 N$5394 VDD p L=2u W=6u
        MN565 N$5394 CK N$5396 GND n L=2u W=6u
        MN571 N$5390 CK N$5392 GND n L=2u W=6u
        MP570 N$5455 CK N$5392 VDD p L=2u W=6u
        MN570 N$5392 N$5391 N$5455 GND n L=2u W=6u
        MN569 N$5397 CK GND GND n L=2u W=6u
        MP569 N$5397 CK VDD VDD p L=2u W=6u
        MN568 N$5393 N$5394 GND GND n L=2u W=6u
        MP568 N$5393 N$5394 VDD VDD p L=2u W=6u
        MN574 N$5388 CK N$5390 GND n L=2u W=6u
        MN573 N$5390 N$5389 GND GND n L=2u W=6u
        MP573 N$5390 N$5389 VDD VDD p L=2u W=6u
        MN572 N$5389 N$5392 GND GND n L=2u W=6u
        MP572 N$5389 N$5392 VDD VDD p L=2u W=6u
        MP571 N$5392 N$5391 N$5390 VDD p L=2u W=6u
        MN577 N$5963 N$5388 GND GND n L=2u W=6u
        MP577 N$5963 N$5388 VDD VDD p L=2u W=6u
        MN576 N$5400 N$5963 GND GND n L=2u W=6u
        MP576 N$5400 N$5963 VDD VDD p L=2u W=6u
        MP607 N$5361 CK N$5363 VDD p L=2u W=6u
        MN607 N$5363 N$5362 N$5361 GND n L=2u W=6u
        MN606 N$5371 CK GND GND n L=2u W=5u
        MP606 N$5371 CK VDD VDD p L=2u W=5u
        MP611 N$5360 N$5362 N$5358 VDD p L=2u W=6u
        MN611 N$5358 CK N$5360 GND n L=2u W=6u
        MN610 N$5360 N$5359 GND GND n L=2u W=6u
        MN583 N$5511 RST GND GND n L=2u W=5u
        MP583 GND N$5385 N$5511 VDD p L=2u W=5u
        MN582 N$5385 RST GND GND n L=2u W=5u
        MN550 N$5408 N$5411 GND GND n L=2u W=6u
        MP550 N$5408 N$5411 VDD VDD p L=2u W=6u
        MP549 N$5411 N$5410 N$5409 VDD p L=2u W=6u
        MN549 N$5409 CK N$5411 GND n L=2u W=6u
        MP555 N$5405 N$5407 VDD VDD p L=2u W=6u
        MN554 N$5406 N$5405 GND GND n L=2u W=6u
        MP554 N$5406 N$5405 VDD VDD p L=2u W=6u
        MP553 N$5407 CK N$5406 VDD p L=2u W=6u
        MN553 N$5406 N$5410 N$5407 GND n L=2u W=6u
        MP552 N$5409 N$5410 N$5407 VDD p L=2u W=6u
        MN557 N$5910 N$5403 GND GND n L=2u W=5u
        MP558 N$5910 N$5963 N$5404 VDD p L=2u W=5u
        MP557 N$5404 N$5403 VDD VDD p L=2u W=5u
        MN556 N$5410 CK GND GND n L=2u W=5u
        MP556 N$5410 CK VDD VDD p L=2u W=5u
        MN555 N$5405 N$5407 GND GND n L=2u W=6u
        MP561 N$5437 CK N$5398 VDD p L=2u W=6u
        MN561 N$5398 N$5397 N$5437 GND n L=2u W=6u
        MN560 N$5399 N$5403 GND GND n L=2u W=5u
        MN559 N$5401 N$5400 N$5399 GND n L=2u W=5u
        MN591 N$5379 N$5387 GND GND n L=2u W=5u
        MP591 N$5379 N$5387 VDD VDD p L=2u W=5u
        MN590 N$5378 N$5379 GND GND n L=2u W=5u
        MP596 N$5381 N$5379 N$5374 VDD p L=2u W=5u
        MN595 N$5375 N$5379 GND GND n L=2u W=5u
        MP595 GND N$5387 N$5375 VDD p L=2u W=5u
        MN594 N$5375 N$5387 N$5413 GND n L=2u W=5u
        MN562 N$5396 CK N$5398 GND n L=2u W=6u
        MN567 N$5403 N$5393 GND GND n L=2u W=6u
        MP567 N$5403 N$5393 VDD VDD p L=2u W=6u
        MP534 N$5423 N$5426 N$5421 VDD p L=2u W=6u
        MN534 N$5421 CK N$5423 GND n L=2u W=6u
        MN533 N$5423 N$5422 GND GND n L=2u W=6u
        MP539 N$5431 CK N$5418 VDD p L=2u W=6u
        MN539 N$5418 N$5417 N$5431 GND n L=2u W=6u
        MN538 N$5426 CK GND GND n L=2u W=5u
        MP538 N$5426 CK VDD VDD p L=2u W=5u
        MN537 N$5419 N$5421 GND GND n L=2u W=6u
        MP537 N$5419 N$5421 VDD VDD p L=2u W=6u
        MN536 N$5420 N$5419 GND GND n L=2u W=6u
        MN542 N$5416 N$5415 GND GND n L=2u W=6u
        MP542 N$5416 N$5415 VDD VDD p L=2u W=6u
        MN541 N$5415 N$5418 GND GND n L=2u W=6u
        MP541 N$5415 N$5418 VDD VDD p L=2u W=6u
        MP540 N$5418 N$5417 N$5416 VDD p L=2u W=6u
        MN540 N$5416 CK N$5418 GND n L=2u W=6u
        MN545 N$5413 N$5412 GND GND n L=2u W=6u
        MP545 N$5413 N$5412 VDD VDD p L=2u W=6u
        MP544 N$5414 CK N$5413 VDD p L=2u W=6u
        MN544 N$5413 N$5417 N$5414 GND n L=2u W=6u
        MP543 N$5416 N$5417 N$5414 VDD p L=2u W=6u
        MP575 N$5388 CK N$5400 VDD p L=2u W=6u
        MN575 N$5400 N$5391 N$5388 GND n L=2u W=6u
        MP574 N$5390 N$5391 N$5388 VDD p L=2u W=6u
        MP580 A5 N$5385 N$5429 VDD p L=2u W=5u
        MN579 N$5387 N$5401 GND GND n L=2u W=6u
        MP579 N$5387 N$5401 VDD VDD p L=2u W=6u
        MN578 N$5391 CK GND GND n L=2u W=5u
        MP578 N$5391 CK VDD VDD p L=2u W=5u
        MN552 N$5407 CK N$5409 GND n L=2u W=6u
        MN551 N$5409 N$5408 GND GND n L=2u W=6u
        MP551 N$5409 N$5408 VDD VDD p L=2u W=6u
        MP520 N$5437 N$5461 N$5438 VDD p L=2u W=6u
        MP519 N$5438 N$5478 N$5439 VDD p L=2u W=6u
        MP518 N$5439 N$5495 N$5442 VDD p L=2u W=6u
        MN523 N$5435 N$5455 GND GND n L=2u W=5u
        MP523 N$5435 N$5455 VDD VDD p L=2u W=5u
        MN522 N$5434 N$5435 N$5475 GND n L=2u W=5u
        MP522 N$5475 N$5455 N$5434 VDD p L=2u W=5u
        MN521 N$5434 N$5455 N$5459 GND n L=2u W=5u
        MP521 N$5459 N$5435 N$5434 VDD p L=2u W=5u
        MN526 N$5431 N$5455 N$5492 GND n L=2u W=5u
        MP526 N$5492 N$5435 N$5431 VDD p L=2u W=5u
        MN525 N$5432 N$5435 N$5492 GND n L=2u W=5u
        MP525 N$5492 N$5455 N$5432 VDD p L=2u W=5u
        MN524 N$5432 N$5455 N$5475 GND n L=2u W=5u
        MP524 N$5475 N$5435 N$5432 VDD p L=2u W=5u
        MN529 N$5430 N$5435 N$5429 GND n L=2u W=5u
        MP529 N$5429 N$5455 N$5430 VDD p L=2u W=5u
        MN528 N$5430 N$5455 N$5511 GND n L=2u W=5u
        MP528 N$5511 N$5435 N$5430 VDD p L=2u W=5u
        MN527 N$5431 N$5435 N$5511 GND n L=2u W=5u
        MP560 N$5401 N$5403 VDD VDD p L=2u W=5u
        MP559 N$5401 N$5400 VDD VDD p L=2u W=5u
        MN558 N$5910 N$5963 GND GND n L=2u W=5u
        MN564 N$5396 N$5395 GND GND n L=2u W=6u
        MP564 N$5396 N$5395 VDD VDD p L=2u W=6u
        MN563 N$5395 N$5398 GND GND n L=2u W=6u
        MP563 N$5395 N$5398 VDD VDD p L=2u W=6u
        MP562 N$5398 N$5397 N$5396 VDD p L=2u W=6u
        MP536 N$5420 N$5419 VDD VDD p L=2u W=6u
        MP535 N$5421 CK N$5420 VDD p L=2u W=6u
        MN535 N$5420 N$5426 N$5421 GND n L=2u W=6u
        MP478 N$5473 N$5474 N$5476 VDD p L=2u W=3u
        MP484 N$5468 N$5474 VDD VDD p L=2u W=3u
        MP483 N$5468 N$5475 VDD VDD p L=2u W=3u
        MP482 N$5468 N$5488 VDD VDD p L=2u W=3u
        MP481 N$5471 N$5472 VDD VDD p L=2u W=3u
        MN481 N$5472 N$5475 N$5469 GND n L=2u W=3u
        MN480 N$5470 N$5474 GND GND n L=2u W=3u
        MN484 N$5464 N$5488 GND GND n L=2u W=3u
        MN483 N$5464 N$5474 GND GND n L=2u W=3u
        MN482 N$5464 N$5475 GND GND n L=2u W=3u
        MP488 N$5465 N$5472 N$5468 VDD p L=2u W=3u
        MP487 N$5465 N$5488 N$5466 VDD p L=2u W=3u
        MP486 N$5466 N$5474 N$5467 VDD p L=2u W=3u
        MP485 N$5467 N$5475 N$5468 VDD p L=2u W=3u
        MN489 N$5461 N$5465 GND GND n L=2u W=3u
        MP489 N$5461 N$5465 VDD VDD p L=2u W=3u
        MN488 N$5465 N$5488 N$5463 GND n L=2u W=3u
        MN487 N$5465 N$5472 N$5464 GND n L=2u W=3u
        MN486 N$5462 N$5474 GND GND n L=2u W=3u
        MN485 N$5463 N$5475 N$5462 GND n L=2u W=3u
        MN490 N$5455 N$5456 GND GND n L=2u W=3u
        MN543 N$5414 CK N$5416 GND n L=2u W=6u
        MP548 N$5434 CK N$5411 VDD p L=2u W=6u
        MN548 N$5411 N$5410 N$5434 GND n L=2u W=6u
        MN547 N$5417 CK GND GND n L=2u W=5u
        MP547 N$5417 CK VDD VDD p L=2u W=5u
        MN546 N$5412 N$5414 GND GND n L=2u W=6u
        MP546 N$5412 N$5414 VDD VDD p L=2u W=6u
        MN519 N$5437 N$5478 GND GND n L=2u W=6u
        MN518 N$5437 N$5495 GND GND n L=2u W=6u
        MN517 N$5437 N$5441 GND GND n L=2u W=6u
        MN49 N$3671 N$3451 GND GND n L=2u W=3u
        MP55 N$3670 N$3664 N$3667 VDD p L=2u W=3u
        MP54 N$3670 GND N$3669 VDD p L=2u W=3u
        MP53 N$3669 N$3701 N$3668 VDD p L=2u W=3u
        MP52 N$3668 N$3451 N$3667 VDD p L=2u W=3u
        MP51 N$3667 N$3701 VDD VDD p L=2u W=3u
        MP50 N$3667 N$3451 VDD VDD p L=2u W=3u
        MP49 N$3667 GND VDD VDD p L=2u W=3u
        MP48 N$3700 N$3664 VDD VDD p L=2u W=3u
        MN48 N$3664 N$3451 N$3666 GND n L=2u W=3u
        MN47 N$3665 N$3701 GND GND n L=2u W=3u
        MN176 N$999 N$995 GND GND n L=2u W=3u
        MN454 N$5498 N$5510 GND GND n L=2u W=3u
        MN453 N$5498 N$5511 GND GND n L=2u W=3u
        MP459 N$5499 N$5508 N$5502 VDD p L=2u W=3u
        MP458 N$5499 N$5507 N$5500 VDD p L=2u W=3u
        MP457 N$5500 N$5510 N$5501 VDD p L=2u W=3u
        MP456 N$5501 N$5511 N$5502 VDD p L=2u W=3u
        MP460 N$5495 N$5499 VDD VDD p L=2u W=3u
        MN459 N$5499 N$5507 N$5497 GND n L=2u W=3u
        MP503 N$5445 N$5449 VDD VDD p L=2u W=3u
        MP517 N$5442 N$5441 N$5440 VDD p L=2u W=6u
        MN507 N$5474 B3 GND GND n L=2u W=3u
        MP507 N$5474 B3 VDD VDD p L=2u W=3u
        MN506 N$5458 GND GND GND n L=2u W=3u
        MP506 N$5458 GND VDD VDD p L=2u W=3u
        MN505 N$5491 B2 GND GND n L=2u W=3u
        MN520 N$5437 N$5461 GND GND n L=2u W=6u
        MN476 N$5471 N$5472 GND GND n L=2u W=3u
        MP480 N$5472 N$5475 N$5473 VDD p L=2u W=3u
        MP479 N$5472 N$5488 N$5476 VDD p L=2u W=3u
        MN57 N$1038 N$6187 N$1041 GND n L=2u W=6u
        MP57 N$1038 N$4988 VDD VDD p L=2u W=6u
        MN141 N$1056 N$4990 GND GND n L=2u W=6u
        MN80 N$2906 N$1035 GND GND n L=2u W=6u
        MP80 N$2906 N$1035 VDD VDD p L=2u W=6u
        MN79 N$1031 N$4989 GND GND n L=2u W=6u
        MN61 N$1044 N$4990 GND GND n L=2u W=6u
        MP61 N$1043 N$6187 VDD VDD p L=2u W=6u
        MN60 N$1043 N$6187 N$1044 GND n L=2u W=6u
        MP60 N$1043 N$4990 VDD VDD p L=2u W=6u
        MN59 N$2905 N$1038 GND GND n L=2u W=6u
        MP59 N$2905 N$1038 VDD VDD p L=2u W=6u
        MN58 N$1041 N$4988 GND GND n L=2u W=6u
        MN64 N$1047 N$4991 GND GND n L=2u W=6u
        MP64 N$1046 N$6187 VDD VDD p L=2u W=6u
        MN63 N$1046 N$6187 N$1047 GND n L=2u W=6u
        MP63 N$1046 N$4991 VDD VDD p L=2u W=6u
        MP3 N$5 N$2907 N$2 VDD p L=2u W=3u
        MP2 N$2 N$2907 VDD VDD p L=2u W=3u
        MP1 N$2 N$4109 VDD VDD p L=2u W=3u
        MP447 N$5512 N$5511 VDD VDD p L=2u W=3u
        MP494 N$5456 N$5459 N$5457 VDD p L=2u W=3u
        MP493 N$5456 N$5471 N$5460 VDD p L=2u W=3u
        MP492 N$5457 N$5458 N$5460 VDD p L=2u W=3u
        MP491 N$5460 N$5458 VDD VDD p L=2u W=3u
        MP490 N$5460 N$5459 VDD VDD p L=2u W=3u
        MP495 N$5455 N$5456 VDD VDD p L=2u W=3u
        MN495 N$5456 N$5459 N$5453 GND n L=2u W=3u
        MN494 N$5454 N$5458 GND GND n L=2u W=3u
        MN52 N$3672 N$3451 N$3673 GND n L=2u W=3u
        MN51 N$3671 GND GND GND n L=2u W=3u
        MN50 N$3671 N$3701 GND GND n L=2u W=3u
        MP282 N$4356 N$4359 VDD VDD p L=2u W=6u
        MN282 N$4356 N$4359 GND GND n L=2u W=6u
        MN283 N$4355 CK N$4356 GND n L=2u W=6u
        MP283 N$4356 N$4360 N$4355 VDD p L=2u W=6u
        MN284 N$4313 N$4360 N$4355 GND n L=2u W=6u
        MP284 N$4355 CK N$4313 VDD p L=2u W=6u
        MP285 N$4313 N$4358 VDD VDD p L=2u W=6u
        MN285 N$4313 N$4358 GND GND n L=2u W=6u
        MP286 N$4358 N$4355 VDD VDD p L=2u W=6u
        MN144 N$1058 N$4991 GND GND n L=2u W=6u
        MN212 N$1067 N$4991 GND GND n L=2u W=6u
        MP144 N$1057 N$5204 VDD VDD p L=2u W=6u
        MN209 N$1065 N$4990 GND GND n L=2u W=6u
        MP209 N$1064 N$5744 VDD VDD p L=2u W=6u
        MN208 N$1064 N$5744 N$1065 GND n L=2u W=6u
        MP208 N$1064 N$4990 VDD VDD p L=2u W=6u
        MN207 N$2902 N$1077 GND GND n L=2u W=6u
        MP167 N$988 N$709 N$987 VDD p L=2u W=3u
        MP28 N$1601 N$31 VDD VDD p L=2u W=3u
        MN34 N$40 N$2904 N$43 GND n L=2u W=3u
        MN33 N$42 N$2906 GND GND n L=2u W=3u
        MN458 N$5499 N$5508 N$5498 GND n L=2u W=3u
        MN457 N$5496 N$5510 GND GND n L=2u W=3u
        MN456 N$5497 N$5511 N$5496 GND n L=2u W=3u
        MN455 N$5498 N$5507 GND GND n L=2u W=3u
        MN461 N$5488 N$5489 GND GND n L=2u W=3u
        MP465 N$5489 N$5492 N$5490 VDD p L=2u W=3u
        MP464 N$5489 N$5505 N$5493 VDD p L=2u W=3u
        MP463 N$5490 N$5491 N$5493 VDD p L=2u W=3u
        MP77 N$2017 N$1034 VDD VDD p L=2u W=6u
        MN76 N$1030 N$4991 GND GND n L=2u W=6u
        MP58 N$1038 N$6187 VDD VDD p L=2u W=6u
        MN154 N$3689 N$1017 N$3692 GND n L=2u W=3u
        MN153 N$3691 N$3456 GND GND n L=2u W=3u
        MN152 N$3692 N$3456 GND GND n L=2u W=3u
        MN151 N$3689 N$3460 N$3691 GND n L=2u W=3u
        MN150 N$3691 N$1017 GND GND n L=2u W=3u
        MN149 N$3690 N$3689 GND GND n L=2u W=3u
        MP153 N$3689 N$1017 N$3688 VDD p L=2u W=3u
        MP454 N$5502 N$5511 VDD VDD p L=2u W=3u
        MN186 N$1011 N$2902 N$1012 GND n L=2u W=3u
        MN185 N$1010 N$2494 GND GND n L=2u W=3u
        MN184 N$1010 N$956 GND GND n L=2u W=3u
        MN190 N$3451 N$1009 GND GND n L=2u W=3u
        MP190 N$3451 N$1009 VDD VDD p L=2u W=3u
        MN165 N$988 N$2903 N$990 GND n L=2u W=3u
        MN189 N$1009 N$2494 N$1011 GND n L=2u W=3u
        MN192 N$1018 N$1607 GND GND n L=2u W=3u
        MN193 N$1016 N$946 N$1018 GND n L=2u W=3u
        MN188 N$1009 N$1002 N$1010 GND n L=2u W=3u
        MN162 N$4321 N$3696 GND GND n L=2u W=3u
        MP162 N$4321 N$3696 VDD VDD p L=2u W=3u
        MP6 N$9 N$6 VDD VDD p L=2u W=3u
        MN6 N$6 N$4109 N$11 GND n L=2u W=3u
        MN5 N$10 N$2907 GND GND n L=2u W=3u
        MN4 N$11 N$2907 GND GND n L=2u W=3u
        MP79 N$1035 N$6186 VDD VDD p L=2u W=6u
        MN78 N$1035 N$6186 N$1031 GND n L=2u W=6u
        MP78 N$1035 N$4989 VDD VDD p L=2u W=6u
        MN77 N$2017 N$1034 GND GND n L=2u W=6u
        MP280 N$4357 N$4360 N$4356 VDD p L=2u W=6u
        MP281 N$4359 N$4357 VDD VDD p L=2u W=6u
        MN281 N$4359 N$4357 GND GND n L=2u W=6u
        MP129 N$3680 N$3700 VDD VDD p L=2u W=3u
        MP128 N$3460 N$3677 VDD VDD p L=2u W=3u
        MN128 N$3677 N$2491 N$3679 GND n L=2u W=3u
        MN127 N$3678 N$3446 GND GND n L=2u W=3u
        MN126 N$3679 N$3446 GND GND n L=2u W=3u
        MN125 N$3677 N$3700 N$3678 GND n L=2u W=3u
        MN124 N$3678 N$2491 GND GND n L=2u W=3u
        MN123 N$3460 N$3677 GND GND n L=2u W=3u
        MP126 N$3677 N$3700 N$3675 VDD p L=2u W=3u
        MN3 N$6 GND N$10 GND n L=2u W=3u
        MN2 N$10 N$4109 GND GND n L=2u W=3u
        MN1 N$9 N$6 GND GND n L=2u W=3u
        MP125 N$3676 N$3446 N$3675 VDD p L=2u W=3u
        MP124 N$3675 N$3446 VDD VDD p L=2u W=3u
        MP123 N$3675 N$2491 VDD VDD p L=2u W=3u
        MN135 N$3683 N$3700 N$3685 GND n L=2u W=3u
        MN56 N$4320 N$3670 GND GND n L=2u W=3u
        MP56 N$4320 N$3670 VDD VDD p L=2u W=3u
        MP127 N$3677 N$2491 N$3676 VDD p L=2u W=3u
        MP117 N$949 N$2908 VDD VDD p L=2u W=3u
        MP118 N$950 N$1579 N$949 VDD p L=2u W=3u
        MN32 N$43 N$2906 GND GND n L=2u W=3u
        MN31 N$40 GND N$42 GND n L=2u W=3u
        MN30 N$42 N$2904 GND GND n L=2u W=3u
        MN29 N$41 N$40 GND GND n L=2u W=3u
        MP33 N$40 N$2904 N$39 VDD p L=2u W=3u
        MP39 N$46 N$2906 N$45 VDD p L=2u W=3u
        MP38 N$45 N$2904 N$44 VDD p L=2u W=3u
        MP37 N$44 N$2906 VDD VDD p L=2u W=3u
        MP156 N$3693 N$1017 VDD VDD p L=2u W=3u
        MP155 N$3693 N$3460 VDD VDD p L=2u W=3u
        MP154 N$3690 N$3689 VDD VDD p L=2u W=3u
        MN243 N$4331 N$4334 N$2020 GND n L=2u W=6u
        MN242 N$4328 CK GND GND n L=2u W=5u
        MP242 N$4328 CK VDD VDD p L=2u W=5u
        MN224 N$4326 N$4323 GND GND n L=2u W=6u
        MP224 N$4326 N$4323 VDD VDD p L=2u W=6u
        MN223 N$4322 N$4326 GND GND n L=2u W=6u
        MP223 N$4322 N$4326 VDD VDD p L=2u W=6u
        MP222 N$4323 CK N$4322 VDD p L=2u W=6u
        MN222 N$4322 N$4328 N$4323 GND n L=2u W=6u
        MN300 N$4368 N$4371 GND GND n L=2u W=6u
        MP300 N$4368 N$4371 VDD VDD p L=2u W=6u
        MN299 N$4371 N$4369 GND GND n L=2u W=6u
        MP299 N$4371 N$4369 VDD VDD p L=2u W=6u
        MP298 N$4369 N$4372 N$4368 VDD p L=2u W=6u
        MN298 N$4368 CK N$4369 GND n L=2u W=6u
        MP297 N$3690 CK N$4369 VDD p L=2u W=6u
        MN297 N$4369 N$4372 N$3690 GND n L=2u W=6u
        MN296 N$4366 CK GND GND n L=2u W=5u
        MP296 N$4366 CK VDD VDD p L=2u W=5u
        MN301 N$4367 CK N$4368 GND n L=2u W=6u
        MN134 N$3683 N$3677 N$3684 GND n L=2u W=3u
        MN161 N$3696 N$3460 N$3698 GND n L=2u W=3u
        MN160 N$3696 N$3689 N$3697 GND n L=2u W=3u
        MN159 N$3699 N$3456 GND GND n L=2u W=3u
        MN158 N$3698 N$1017 N$3699 GND n L=2u W=3u
        MN157 N$3697 N$3460 GND GND n L=2u W=3u
        MN156 N$3697 N$3456 GND GND n L=2u W=3u
        MN155 N$3697 N$1017 GND GND n L=2u W=3u
        MN187 N$1012 N$956 GND GND n L=2u W=3u
        MP132 N$3681 N$2491 N$3680 VDD p L=2u W=3u
        MP131 N$3680 N$3446 VDD VDD p L=2u W=3u
        MP130 N$3680 N$2491 VDD VDD p L=2u W=3u
        MN104 N$940 N$1578 N$941 GND n L=2u W=3u
        MN148 N$1584 N$1059 GND GND n L=2u W=6u
        MP148 N$1584 N$1059 VDD VDD p L=2u W=6u
        MN147 N$1060 N$4989 GND GND n L=2u W=6u
        MP147 N$1059 N$5204 VDD VDD p L=2u W=6u
        MN146 N$1059 N$5204 N$1060 GND n L=2u W=6u
        MP146 N$1059 N$4989 VDD VDD p L=2u W=6u
        MN145 N$1579 N$1057 GND GND n L=2u W=6u
        MP145 N$1579 N$1057 VDD VDD p L=2u W=6u
        MP455 N$5502 N$5510 VDD VDD p L=2u W=3u
        MN137 N$1051 N$5204 N$1053 GND n L=2u W=6u
        MP137 N$1051 N$4988 VDD VDD p L=2u W=6u
        MP139 N$1578 N$1051 VDD VDD p L=2u W=6u
        MN138 N$1053 N$4988 GND GND n L=2u W=6u
        MP71 N$2907 N$1033 VDD VDD p L=2u W=6u
        MN70 N$1029 N$4988 GND GND n L=2u W=6u
        MP70 N$1033 N$6186 VDD VDD p L=2u W=6u
        MN69 N$1033 N$6186 N$1029 GND n L=2u W=6u
        MP69 N$1033 N$4988 VDD VDD p L=2u W=6u
        MN143 N$1057 N$5204 N$1058 GND n L=2u W=6u
        MP213 N$1607 N$1066 VDD VDD p L=2u W=6u
        MN73 N$1028 N$4990 GND GND n L=2u W=6u
        MN13 N$15 GND N$17 GND n L=2u W=3u
        MN12 N$15 N$6 N$16 GND n L=2u W=3u
        MN11 N$18 N$2907 GND GND n L=2u W=3u
        MP116 N$949 N$1579 VDD VDD p L=2u W=3u
        MP5 N$6 N$4109 N$5 VDD p L=2u W=3u
        MP4 N$6 GND N$2 VDD p L=2u W=3u
        MP157 N$3693 N$3456 VDD VDD p L=2u W=3u
        MP244 N$4331 N$4334 N$4330 VDD p L=2u W=6u
        MN244 N$4330 CK N$4331 GND n L=2u W=6u
        MP243 N$2020 CK N$4331 VDD p L=2u W=6u
        MP141 N$1055 N$5204 VDD VDD p L=2u W=6u
        MN140 N$1055 N$5204 N$1056 GND n L=2u W=6u
        MP140 N$1055 N$4990 VDD VDD p L=2u W=6u
        MN139 N$1578 N$1051 GND GND n L=2u W=6u
        MP86 N$2903 N$916 VDD VDD p L=2u W=3u
        MN86 N$916 N$707 N$920 GND n L=2u W=3u
        MP87 N$921 N$9 VDD VDD p L=2u W=3u
        MP88 N$921 N$707 VDD VDD p L=2u W=3u
        MP89 N$921 N$1601 VDD VDD p L=2u W=3u
        MP90 N$922 N$707 N$921 VDD p L=2u W=3u
        MN195 N$1018 N$1584 GND GND n L=2u W=3u
        MN194 N$1019 N$1584 GND GND n L=2u W=3u
        MN197 N$1024 N$1607 GND GND n L=2u W=3u
        MP203 N$1023 N$1016 N$1020 VDD p L=2u W=3u
        MP202 N$1023 N$946 N$1022 VDD p L=2u W=3u
        MP201 N$1022 N$1584 N$1021 VDD p L=2u W=3u
        MP200 N$1021 N$1607 N$1020 VDD p L=2u W=3u
        MP199 N$1020 N$1584 VDD VDD p L=2u W=3u
        MN203 N$1023 N$946 N$1025 GND n L=2u W=3u
        MN202 N$1023 N$1016 N$1024 GND n L=2u W=3u
        MN201 N$1026 N$1584 GND GND n L=2u W=3u
        MN133 N$3686 N$3446 GND GND n L=2u W=3u
        MN132 N$3685 N$2491 N$3686 GND n L=2u W=3u
        MN131 N$3684 N$3700 GND GND n L=2u W=3u
        MN130 N$3684 N$3446 GND GND n L=2u W=3u
        MN129 N$3684 N$2491 GND GND n L=2u W=3u
        MP135 N$3683 N$3677 N$3680 VDD p L=2u W=3u
        MP134 N$3683 N$3700 N$3682 VDD p L=2u W=3u
        MP133 N$3682 N$3446 N$3681 VDD p L=2u W=3u
        MP206 N$1077 N$5744 VDD VDD p L=2u W=6u
        MN205 N$1077 N$5744 N$1062 GND n L=2u W=6u
        MP205 N$1077 N$4988 VDD VDD p L=2u W=6u
        MP31 N$39 N$2906 N$36 VDD p L=2u W=3u
        MP165 N$987 N$942 N$986 VDD p L=2u W=3u
        MP164 N$986 N$942 VDD VDD p L=2u W=3u
        MP163 N$986 N$709 VDD VDD p L=2u W=3u
        MN39 N$50 N$2906 GND GND n L=2u W=3u
        MP207 N$2902 N$1077 VDD VDD p L=2u W=6u
        MP8 N$12 N$4109 VDD VDD p L=2u W=3u
        MP11 N$14 N$2907 N$13 VDD p L=2u W=3u
        MP7 N$12 GND VDD VDD p L=2u W=3u
        MN8 N$16 N$2907 GND GND n L=2u W=3u
        MN181 N$1004 N$956 GND GND n L=2u W=3u
        MN180 N$1005 N$956 GND GND n L=2u W=3u
        MN179 N$1002 N$2494 N$1004 GND n L=2u W=3u
        MN178 N$1004 N$2902 GND GND n L=2u W=3u
        MN177 N$3446 N$1002 GND GND n L=2u W=3u
        MP166 N$988 N$2903 N$986 VDD p L=2u W=3u
        MN191 N$1017 N$1016 GND GND n L=2u W=3u
        MP181 N$1002 N$2902 N$1001 VDD p L=2u W=3u
        MP180 N$1002 N$2494 N$1000 VDD p L=2u W=3u
        MP179 N$1001 N$956 N$1000 VDD p L=2u W=3u
        MP178 N$1000 N$956 VDD VDD p L=2u W=3u
        MN216 N$3456 N$1068 GND GND n L=2u W=6u
        MP216 N$3456 N$1068 VDD VDD p L=2u W=6u
        MP247 N$4330 N$4334 N$4329 VDD p L=2u W=6u
        MN247 N$4329 CK N$4330 GND n L=2u W=6u
        MN246 N$4330 N$4333 GND GND n L=2u W=6u
        MP246 N$4330 N$4333 VDD VDD p L=2u W=6u
        MN245 N$4333 N$4331 GND GND n L=2u W=6u
        MP245 N$4333 N$4331 VDD VDD p L=2u W=6u
        MN107 N$938 N$25 N$940 GND n L=2u W=3u
        MN106 N$938 N$932 N$939 GND n L=2u W=3u
        MN105 N$941 N$51 GND GND n L=2u W=3u
        MP29 N$36 N$2904 VDD VDD p L=2u W=3u
        MP30 N$36 N$2906 VDD VDD p L=2u W=3u
        MP103 N$935 N$51 VDD VDD p L=2u W=3u
        MP102 N$935 N$1578 VDD VDD p L=2u W=3u
        MP101 N$935 N$25 VDD VDD p L=2u W=3u
        MP100 N$2494 N$932 VDD VDD p L=2u W=3u
        MN100 N$932 N$1578 N$934 GND n L=2u W=3u
        MN99 N$933 N$51 GND GND n L=2u W=3u
        MN98 N$934 N$51 GND GND n L=2u W=3u
        MN97 N$932 N$25 N$933 GND n L=2u W=3u
        MP184 N$1006 N$2902 VDD VDD p L=2u W=3u
        MP183 N$1006 N$2494 VDD VDD p L=2u W=3u
        MP182 N$3446 N$1002 VDD VDD p L=2u W=3u
        MN204 N$2491 N$1023 GND GND n L=2u W=3u
        MP204 N$2491 N$1023 VDD VDD p L=2u W=3u
        MN182 N$1002 N$2902 N$1005 GND n L=2u W=3u
        MN85 N$919 N$1601 GND GND n L=2u W=3u
        MN84 N$920 N$1601 GND GND n L=2u W=3u
        MN83 N$916 N$9 N$919 GND n L=2u W=3u
        MN82 N$919 N$707 GND GND n L=2u W=3u
        MN81 N$2903 N$916 GND GND n L=2u W=3u
        MN200 N$1025 N$1607 N$1026 GND n L=2u W=3u
        MN199 N$1024 N$946 GND GND n L=2u W=3u
        MN198 N$1024 N$1584 GND GND n L=2u W=3u
        MN103 N$939 N$25 GND GND n L=2u W=3u
        MN102 N$939 N$51 GND GND n L=2u W=3u
        MN101 N$939 N$1578 GND GND n L=2u W=3u
        MN196 N$1016 N$1607 N$1019 GND n L=2u W=3u
        MN206 N$1062 N$4988 GND GND n L=2u W=6u
        MN90 N$926 N$707 N$927 GND n L=2u W=3u
        MP104 N$936 N$1578 N$935 VDD p L=2u W=3u
        MP32 N$40 GND N$36 VDD p L=2u W=3u
        MP21 N$28 GND VDD VDD p L=2u W=3u
        MP20 N$25 N$24 VDD VDD p L=2u W=3u
        MN20 N$24 N$2905 N$27 GND n L=2u W=3u
        MN19 N$26 N$2017 GND GND n L=2u W=3u
        MN18 N$27 N$2017 GND GND n L=2u W=3u
        MN17 N$24 GND N$26 GND n L=2u W=3u
        MP27 N$31 N$24 N$28 VDD p L=2u W=3u
        MP26 N$31 GND N$30 VDD p L=2u W=3u
        MP25 N$30 N$2017 N$29 VDD p L=2u W=3u
        MP24 N$29 N$2905 N$28 VDD p L=2u W=3u
        MN7 N$16 N$4109 GND GND n L=2u W=3u
        MP13 N$15 N$6 N$12 VDD p L=2u W=3u
        MP12 N$15 GND N$14 VDD p L=2u W=3u
        MN9 N$16 GND GND GND n L=2u W=3u
        MN10 N$17 N$4109 N$18 GND n L=2u W=3u
        MP10 N$13 N$4109 N$12 VDD p L=2u W=3u
        MP9 N$12 N$2907 VDD VDD p L=2u W=3u
        MN41 N$47 GND N$49 GND n L=2u W=3u
        MN40 N$47 N$40 N$48 GND n L=2u W=3u
        MP42 N$51 N$47 VDD VDD p L=2u W=3u
        MN42 N$51 N$47 GND GND n L=2u W=3u
        MP177 N$1000 N$2902 VDD VDD p L=2u W=3u
        MN163 N$3701 N$988 GND GND n L=2u W=3u
        MN164 N$990 N$709 GND GND n L=2u W=3u
        MN167 N$990 N$942 GND GND n L=2u W=3u
        MN166 N$991 N$942 GND GND n L=2u W=3u
        MN170 N$996 N$942 GND GND n L=2u W=3u
        MN169 N$996 N$709 GND GND n L=2u W=3u
        MP175 N$995 N$988 N$992 VDD p L=2u W=3u
        MN210 N$709 N$1064 GND GND n L=2u W=6u
        MP210 N$709 N$1064 VDD VDD p L=2u W=6u
        MN28 N$1601 N$31 GND GND n L=2u W=3u
        MN88 N$925 N$1601 GND GND n L=2u W=3u
        MN87 N$925 N$707 GND GND n L=2u W=3u
        MP93 N$924 N$916 N$921 VDD p L=2u W=3u
        MP92 N$924 N$9 N$923 VDD p L=2u W=3u
        MP91 N$923 N$1601 N$922 VDD p L=2u W=3u
        MP161 N$3696 N$3689 N$3693 VDD p L=2u W=3u
        MP160 N$3696 N$3460 N$3695 VDD p L=2u W=3u
        MP159 N$3695 N$3456 N$3694 VDD p L=2u W=3u
        MP158 N$3694 N$1017 N$3693 VDD p L=2u W=3u
        MN68 N$2908 N$1049 GND GND n L=2u W=6u
        MP23 N$28 N$2017 VDD VDD p L=2u W=3u
        MP22 N$28 N$2905 VDD VDD p L=2u W=3u
        MN27 N$31 GND N$33 GND n L=2u W=3u
        MN26 N$31 N$24 N$32 GND n L=2u W=3u
        MN25 N$34 N$2017 GND GND n L=2u W=3u
        MN24 N$33 N$2905 N$34 GND n L=2u W=3u
        MN23 N$32 GND GND GND n L=2u W=3u
        MN22 N$32 N$2017 GND GND n L=2u W=3u
        MP107 N$938 N$932 N$935 VDD p L=2u W=3u
        MP106 N$938 N$25 N$937 VDD p L=2u W=3u
        MP105 N$937 N$51 N$936 VDD p L=2u W=3u
        MP85 N$916 N$707 N$915 VDD p L=2u W=3u
        MP84 N$916 N$9 N$914 VDD p L=2u W=3u
        MP83 N$915 N$1601 N$914 VDD p L=2u W=3u
        MN118 N$954 N$1579 N$955 GND n L=2u W=3u
        MN117 N$953 N$41 GND GND n L=2u W=3u
        MN93 N$924 N$9 N$926 GND n L=2u W=3u
        MN92 N$924 N$916 N$925 GND n L=2u W=3u
        MN91 N$927 N$1601 GND GND n L=2u W=3u
        MP17 N$23 N$2017 N$20 VDD p L=2u W=3u
        MP16 N$20 N$2017 VDD VDD p L=2u W=3u
        MP15 N$20 N$2905 VDD VDD p L=2u W=3u
        MP259 N$4338 N$4335 VDD VDD p L=2u W=6u
        MN258 N$4312 N$4338 GND GND n L=2u W=6u
        MP258 N$4312 N$4338 VDD VDD p L=2u W=6u
        MP257 N$4335 CK N$4312 VDD p L=2u W=6u
        MN257 N$4312 N$4340 N$4335 GND n L=2u W=6u
        MP256 N$4336 N$4340 N$4335 VDD p L=2u W=6u
        MN256 N$4335 CK N$4336 GND n L=2u W=6u
        MN255 N$4336 N$4339 GND GND n L=2u W=6u
        MP255 N$4336 N$4339 VDD VDD p L=2u W=6u
        MN254 N$4339 N$4337 GND GND n L=2u W=6u
        MP221 N$4324 N$4328 N$4323 VDD p L=2u W=6u
        MN221 N$4323 CK N$4324 GND n L=2u W=6u
        MN220 N$4324 N$4327 GND GND n L=2u W=6u
        MP220 N$4324 N$4327 VDD VDD p L=2u W=6u
        MN219 N$4327 N$4325 GND GND n L=2u W=6u
        MP219 N$4327 N$4325 VDD VDD p L=2u W=6u
        MP218 N$4325 N$4328 N$4324 VDD p L=2u W=6u
        MN218 N$4324 CK N$4325 GND n L=2u W=6u
        MP217 N$37 CK N$4325 VDD p L=2u W=6u
        MN217 N$4325 N$4328 N$37 GND n L=2u W=6u
        MP143 N$1057 N$4991 VDD VDD p L=2u W=6u
        MP169 N$992 N$2903 VDD VDD p L=2u W=3u
        MP168 N$3701 N$988 VDD VDD p L=2u W=3u
        MN168 N$988 N$709 N$991 GND n L=2u W=3u
        MP40 N$47 GND N$46 VDD p L=2u W=3u
        MN21 N$32 N$2905 GND GND n L=2u W=3u
        MP212 N$1066 N$5744 VDD VDD p L=2u W=6u
        MN211 N$1066 N$5744 N$1067 GND n L=2u W=6u
        MP211 N$1066 N$4991 VDD VDD p L=2u W=6u
        MP66 N$1049 N$4989 VDD VDD p L=2u W=6u
        MN65 N$2904 N$1046 GND GND n L=2u W=6u
        MP65 N$2904 N$1046 VDD VDD p L=2u W=6u
        MP291 N$4362 N$4365 VDD VDD p L=2u W=6u
        MN290 N$4365 N$4363 GND GND n L=2u W=6u
        MP290 N$4365 N$4363 VDD VDD p L=2u W=6u
        MP289 N$4363 N$4366 N$4362 VDD p L=2u W=6u
        MN289 N$4362 CK N$4363 GND n L=2u W=6u
        MP288 N$4321 CK N$4363 VDD p L=2u W=6u
        MN288 N$4363 N$4366 N$4321 GND n L=2u W=6u
        MN287 N$4360 CK GND GND n L=2u W=5u
        MP287 N$4360 CK VDD VDD p L=2u W=5u
        MN286 N$4358 N$4355 GND GND n L=2u W=6u
        MP254 N$4339 N$4337 VDD VDD p L=2u W=6u
        MP253 N$4337 N$4340 N$4336 VDD p L=2u W=6u
        MN253 N$4336 CK N$4337 GND n L=2u W=6u
        MP252 N$928 CK N$4337 VDD p L=2u W=6u
        MN252 N$4337 N$4340 N$928 GND n L=2u W=6u
        MN251 N$4334 CK GND GND n L=2u W=5u
        MP251 N$4334 CK VDD VDD p L=2u W=5u
        MN250 N$4332 N$4329 GND GND n L=2u W=6u
        MP250 N$4332 N$4329 VDD VDD p L=2u W=6u
        MN249 N$4311 N$4332 GND GND n L=2u W=6u
        MP249 N$4311 N$4332 VDD VDD p L=2u W=6u
        MP198 N$1020 N$1607 VDD VDD p L=2u W=3u
        MP197 N$1020 N$946 VDD VDD p L=2u W=3u
        MP196 N$1017 N$1016 VDD VDD p L=2u W=3u
        MN94 N$928 N$924 GND GND n L=2u W=3u
        MP94 N$928 N$924 VDD VDD p L=2u W=3u
        MN14 N$2020 N$15 GND GND n L=2u W=3u
        MP14 N$2020 N$15 VDD VDD p L=2u W=3u
        MP119 N$951 N$2908 N$950 VDD p L=2u W=3u
        MN260 N$4340 CK GND GND n L=2u W=5u
        MP260 N$4340 CK VDD VDD p L=2u W=5u
        MN259 N$4338 N$4335 GND GND n L=2u W=6u
        MP407 N$5927 N$5932 N$5934 VDD p L=2u W=5u
        MN406 N$5934 N$5932 N$5925 GND n L=2u W=5u
        MP406 N$5925 N$5349 N$5934 VDD p L=2u W=5u
        MN369 N$5933 N$5349 N$5926 GND n L=2u W=5u
        MP369 N$5926 N$5932 N$5933 VDD p L=2u W=5u
        MN368 N$5933 N$5932 N$5924 GND n L=2u W=5u
        MP368 N$5924 N$5349 N$5933 VDD p L=2u W=5u
        MN367 N$5932 N$5349 GND GND n L=2u W=5u
        MP367 N$5932 N$5349 VDD VDD p L=2u W=5u
        MN366 N$5931 N$5349 N$5925 GND n L=2u W=5u
        MP366 N$5925 N$5932 N$5931 VDD p L=2u W=5u
        MN365 N$5931 N$5932 N$5922 GND n L=2u W=5u
        MP365 N$5922 N$5349 N$5931 VDD p L=2u W=5u
        MN364 N$5930 N$5357 GND GND n L=2u W=5u
        MP364 GND N$5923 N$5930 VDD p L=2u W=5u
        MN363 N$5930 N$5923 N$5920 GND n L=2u W=5u
        MP363 N$5920 N$5357 N$5930 VDD p L=2u W=5u
        MN362 N$5929 N$5357 N$5920 GND n L=2u W=5u
        MP362 N$5920 N$5923 N$5929 VDD p L=2u W=5u
        MN361 N$5929 N$5923 N$5919 GND n L=2u W=5u
        MP361 N$5919 N$5357 N$5929 VDD p L=2u W=5u
        MP114 N$946 N$945 VDD VDD p L=2u W=3u
        MP115 N$949 N$41 VDD VDD p L=2u W=3u
        MN263 N$4346 N$4344 GND GND n L=2u W=6u
        MP263 N$4346 N$4344 VDD VDD p L=2u W=6u
        MP262 N$4344 N$4347 N$4343 VDD p L=2u W=6u
        MN262 N$4343 CK N$4344 GND n L=2u W=6u
        MP261 N$999 CK N$4344 VDD p L=2u W=6u
        MN261 N$4344 N$4347 N$999 GND n L=2u W=6u
        MP292 N$4362 N$4366 N$4361 VDD p L=2u W=6u
        MN292 N$4361 CK N$4362 GND n L=2u W=6u
        MN291 N$4362 N$4365 GND GND n L=2u W=6u
        MP423 N$5934 N$5341 N$5897 VDD p L=2u W=5u
        MN422 N$5942 N$5341 N$5936 GND n L=2u W=5u
        MP422 N$5936 N$5941 N$5942 VDD p L=2u W=5u
        MN421 N$5942 N$5941 N$5933 GND n L=2u W=5u
        MP421 N$5933 N$5341 N$5942 VDD p L=2u W=5u
        MN420 N$5941 N$5341 GND GND n L=2u W=5u
        MP420 N$5941 N$5341 VDD VDD p L=2u W=5u
        MN419 N$5956 N$5341 N$5935 GND n L=2u W=5u
        MP419 N$5935 N$5941 N$5956 VDD p L=2u W=5u
        MN418 N$5956 N$5941 N$5931 GND n L=2u W=5u
        MP418 N$5931 N$5341 N$5956 VDD p L=2u W=5u
        MN417 N$5939 N$5349 GND GND n L=2u W=5u
        MP417 GND N$5932 N$5939 VDD p L=2u W=5u
        MN416 N$5939 N$5932 N$5930 GND n L=2u W=5u
        MP416 N$5930 N$5349 N$5939 VDD p L=2u W=5u
        MN415 N$5938 N$5349 GND GND n L=2u W=5u
        MP415 GND N$5932 N$5938 VDD p L=2u W=5u
        MN414 N$5938 N$5932 N$5929 GND n L=2u W=5u
        MP414 N$5929 N$5349 N$5938 VDD p L=2u W=5u
        MN413 N$5937 N$5349 N$5930 GND n L=2u W=5u
        MP413 N$5930 N$5932 N$5937 VDD p L=2u W=5u
        MP248 N$4329 CK N$4311 VDD p L=2u W=6u
        MN248 N$4311 N$4334 N$4329 GND n L=2u W=6u
        MP279 N$3704 CK N$4357 VDD p L=2u W=6u
        MN279 N$4357 N$4360 N$3704 GND n L=2u W=6u
        MN278 N$4354 CK GND GND n L=2u W=5u
        MP278 N$4354 CK VDD VDD p L=2u W=5u
        MN277 N$4352 N$4349 GND GND n L=2u W=6u
        MP277 N$4352 N$4349 VDD VDD p L=2u W=6u
        MN408 N$5935 N$5932 N$5926 GND n L=2u W=5u
        MP408 N$5926 N$5349 N$5935 VDD p L=2u W=5u
        MN407 N$5934 N$5349 N$5927 GND n L=2u W=5u
        MN269 N$4347 CK GND GND n L=2u W=5u
        MP269 N$4347 CK VDD VDD p L=2u W=5u
        MN268 N$4345 N$4342 GND GND n L=2u W=6u
        MP268 N$4345 N$4342 VDD VDD p L=2u W=6u
        MN267 N$4341 N$4345 GND GND n L=2u W=6u
        MP267 N$4341 N$4345 VDD VDD p L=2u W=6u
        MP266 N$4342 CK N$4341 VDD p L=2u W=6u
        MN266 N$4341 N$4347 N$4342 GND n L=2u W=6u
        MP265 N$4343 N$4347 N$4342 VDD p L=2u W=6u
        MN265 N$4342 CK N$4343 GND n L=2u W=6u
        MN264 N$4343 N$4346 GND GND n L=2u W=6u
        MP264 N$4343 N$4346 VDD VDD p L=2u W=6u
        MN295 N$4364 N$4361 GND GND n L=2u W=6u
        MP295 N$4364 N$4361 VDD VDD p L=2u W=6u
        MN294 N$4314 N$4364 GND GND n L=2u W=6u
        MP294 N$4314 N$4364 VDD VDD p L=2u W=6u
        MP293 N$4361 CK N$4314 VDD p L=2u W=6u
        MN293 N$4314 N$4366 N$4361 GND n L=2u W=6u
        MP381 N$5765 N$5948 N$5764 VDD p L=2u W=3u
        MP380 N$5764 N$5948 VDD VDD p L=2u W=3u
        MN434 N$5948 N$5341 GND GND n L=2u W=5u
        MP634 N$5420 N$5338 N$5337 VDD p L=2u W=5u
        MN639 N$5334 N$5910 N$5381 GND n L=2u W=5u
        MP639 N$5381 N$5338 N$5334 VDD p L=2u W=5u
        MN638 N$5335 N$5338 GND GND n L=2u W=5u
        MP638 GND N$5910 N$5335 VDD p L=2u W=5u
        MN637 N$5335 N$5910 N$5413 GND n L=2u W=5u
        MP637 N$5413 N$5338 N$5335 VDD p L=2u W=5u
        MN471 N$5479 N$5491 GND GND n L=2u W=3u
        MP461 N$5493 N$5492 VDD VDD p L=2u W=3u
        MN460 N$5495 N$5499 GND GND n L=2u W=3u
        MN393 N$5785 N$5783 GND GND n L=2u W=3u
        MP397 N$5783 N$4311 N$5782 VDD p L=2u W=3u
        MP396 N$5783 N$5769 N$5781 VDD p L=2u W=3u
        MP395 N$5782 N$5951 N$5781 VDD p L=2u W=3u
        MP394 N$5781 N$5951 VDD VDD p L=2u W=3u
        MP401 N$5788 N$5951 VDD VDD p L=2u W=3u
        MP400 N$5788 N$4311 VDD VDD p L=2u W=3u
        MP399 N$5788 N$5769 VDD VDD p L=2u W=3u
        MP398 N$5785 N$5783 VDD VDD p L=2u W=3u
        MN398 N$5783 N$4311 N$5787 GND n L=2u W=3u
        MN397 N$5786 N$5951 GND GND n L=2u W=3u
        MN396 N$5787 N$5951 GND GND n L=2u W=3u
        MN400 N$5792 N$5951 GND GND n L=2u W=3u
        MN399 N$5792 N$4311 GND GND n L=2u W=3u
        MP405 N$5791 N$5783 N$5788 VDD p L=2u W=3u
        MP404 N$5791 N$5769 N$5790 VDD p L=2u W=3u
        MP403 N$5790 N$5951 N$5789 VDD p L=2u W=3u
        MP402 N$5789 N$4311 N$5788 VDD p L=2u W=3u
        MP474 OUT1 N$5791 VDD VDD p L=2u W=3u
        MN405 N$5791 N$5769 N$5793 GND n L=2u W=3u
        MN475 N$5478 N$5482 GND GND n L=2u W=3u
        MP475 N$5478 N$5482 VDD VDD p L=2u W=3u
        MN473 N$5482 N$5505 N$5480 GND n L=2u W=3u
        MN479 N$5469 N$5474 GND GND n L=2u W=3u
        MN478 N$5472 N$5488 N$5470 GND n L=2u W=3u
        MN477 N$5470 N$5475 GND GND n L=2u W=3u
        MP383 N$5766 N$4322 N$5765 VDD p L=2u W=3u
        MP382 N$5766 GND N$5764 VDD p L=2u W=3u
        MN270 N$4351 N$4354 N$4320 GND n L=2u W=6u
        MP513 N$5801 N$5799 VDD VDD p L=2u W=3u
        MN513 N$5799 N$4312 N$5803 GND n L=2u W=3u
        MN512 N$5802 N$5945 GND GND n L=2u W=3u
        MN511 N$5803 N$5945 GND GND n L=2u W=3u
        MN510 N$5799 N$5785 N$5802 GND n L=2u W=3u
        MN509 N$5802 N$4312 GND GND n L=2u W=3u
        MN508 N$5801 N$5799 GND GND n L=2u W=3u
        MP776 N$5807 N$5785 N$5806 VDD p L=2u W=3u
        MP775 N$5806 N$5945 N$5805 VDD p L=2u W=3u
        MP774 N$5805 N$4312 N$5804 VDD p L=2u W=3u
        MP516 N$5804 N$5945 VDD VDD p L=2u W=3u
        MP515 N$5804 N$4312 VDD VDD p L=2u W=3u
        MP514 N$5804 N$5785 VDD VDD p L=2u W=3u
        MN775 N$5810 N$5945 GND GND n L=2u W=3u
        MN774 N$5809 N$4312 N$5810 GND n L=2u W=3u
        MN516 N$5808 N$5785 GND GND n L=2u W=3u
        MN515 N$5808 N$5945 GND GND n L=2u W=3u
        MN514 N$5808 N$4312 GND GND n L=2u W=3u
        MP777 N$5807 N$5799 N$5804 VDD p L=2u W=3u
        MP780 N$5813 N$5955 VDD VDD p L=2u W=3u
        MP779 N$5813 N$4341 VDD VDD p L=2u W=3u
        MN385 N$5776 N$4322 GND GND n L=2u W=3u
        MP391 N$5775 N$5766 N$5772 VDD p L=2u W=3u
        MP393 N$5781 N$4311 VDD VDD p L=2u W=3u
        MN392 OUT0 N$5775 GND GND n L=2u W=3u
        MP392 OUT0 N$5775 VDD VDD p L=2u W=3u
        MN391 N$5775 GND N$5777 GND n L=2u W=3u
        MN390 N$5775 N$5766 N$5776 GND n L=2u W=3u
        MN395 N$5783 N$5769 N$5786 GND n L=2u W=3u
        MN394 N$5786 N$4311 GND GND n L=2u W=3u
        MP781 N$5814 N$5955 N$5813 VDD p L=2u W=3u
        MP787 N$5820 N$5955 VDD VDD p L=2u W=3u
        MP786 N$5820 N$4341 VDD VDD p L=2u W=3u
        MP785 N$5820 N$5801 VDD VDD p L=2u W=3u
        MP784 N$5817 N$5815 VDD VDD p L=2u W=3u
        MN784 N$5815 N$4341 N$5819 GND n L=2u W=3u
        MN783 N$5818 N$5955 GND GND n L=2u W=3u
        MN782 N$5819 N$5955 GND GND n L=2u W=3u
        MN786 N$5824 N$5955 GND GND n L=2u W=3u
        MN785 N$5824 N$4341 GND GND n L=2u W=3u
        MP791 N$5823 N$5815 N$5820 VDD p L=2u W=3u
        MP790 N$5823 N$5801 N$5822 VDD p L=2u W=3u
        MP789 N$5822 N$5955 N$5821 VDD p L=2u W=3u
        MP788 N$5821 N$4341 N$5820 VDD p L=2u W=3u
        MN792 OUT3 N$5823 GND GND n L=2u W=3u
        MP792 OUT3 N$5823 VDD VDD p L=2u W=3u
        MN791 N$5823 N$5801 N$5825 GND n L=2u W=3u
        MN790 N$5823 N$5815 N$5824 GND n L=2u W=3u
        MN789 N$5826 N$5955 GND GND n L=2u W=3u
        MN788 N$5825 N$4341 N$5826 GND n L=2u W=3u
        MN787 N$5824 N$5801 GND GND n L=2u W=3u
        MN404 N$5791 N$5783 N$5792 GND n L=2u W=3u
        MN403 N$5794 N$5951 GND GND n L=2u W=3u
        MN402 N$5793 N$4311 N$5794 GND n L=2u W=3u
        MN401 N$5792 N$5769 GND GND n L=2u W=3u
        MP512 N$5799 N$4312 N$5798 VDD p L=2u W=3u
        MP511 N$5799 N$5785 N$5797 VDD p L=2u W=3u
        MP510 N$5798 N$5945 N$5797 VDD p L=2u W=3u
        MP509 N$5797 N$5945 VDD VDD p L=2u W=3u
        MP508 N$5797 N$4312 VDD VDD p L=2u W=3u
        MN474 OUT1 N$5791 GND GND n L=2u W=3u
        MN795 N$5831 N$5817 N$5834 GND n L=2u W=3u
        MN794 N$5834 N$4348 GND GND n L=2u W=3u
        MN793 N$5833 N$5831 GND GND n L=2u W=3u
        MP803 N$5838 N$5896 N$5837 VDD p L=2u W=3u
        MP802 N$5837 N$4348 N$5836 VDD p L=2u W=3u
        MP801 N$5836 N$5896 VDD VDD p L=2u W=3u
        MP800 N$5836 N$4348 VDD VDD p L=2u W=3u
        MP799 N$5836 N$5817 VDD VDD p L=2u W=3u
        MN803 N$5842 N$5896 GND GND n L=2u W=3u
        MN802 N$5841 N$4348 N$5842 GND n L=2u W=3u
        MN801 N$5840 N$5817 GND GND n L=2u W=3u
        MN800 N$5840 N$5896 GND GND n L=2u W=3u
        MN799 N$5840 N$4348 GND GND n L=2u W=3u
        MP805 N$5839 N$5831 N$5836 VDD p L=2u W=3u
        MP804 N$5839 N$5817 N$5838 VDD p L=2u W=3u
        MP808 N$5845 N$5897 VDD VDD p L=2u W=3u
        MP807 N$5845 N$4313 VDD VDD p L=2u W=3u
        MN806 OUT4 N$5839 GND GND n L=2u W=3u
        MP806 OUT4 N$5839 VDD VDD p L=2u W=3u
        MN778 OUT2 N$5807 GND GND n L=2u W=3u
        MP778 OUT2 N$5807 VDD VDD p L=2u W=3u
        MN777 N$5807 N$5785 N$5809 GND n L=2u W=3u
        MN776 N$5807 N$5799 N$5808 GND n L=2u W=3u
        MN781 N$5815 N$5801 N$5818 GND n L=2u W=3u
        MN780 N$5818 N$4341 GND GND n L=2u W=3u
        MN779 N$5817 N$5815 GND GND n L=2u W=3u
        MP783 N$5815 N$4341 N$5814 VDD p L=2u W=3u
        MP782 N$5815 N$5801 N$5813 VDD p L=2u W=3u
        MP812 N$5849 N$5847 VDD VDD p L=2u W=3u
        MN812 N$5847 N$4313 N$5851 GND n L=2u W=3u
        MN811 N$5850 N$5897 GND GND n L=2u W=3u
        MN810 N$5851 N$5897 GND GND n L=2u W=3u
        MN814 N$5856 N$5897 GND GND n L=2u W=3u
        MN813 N$5856 N$4313 GND GND n L=2u W=3u
        MP819 N$5855 N$5847 N$5852 VDD p L=2u W=3u
        MP818 N$5855 N$5833 N$5854 VDD p L=2u W=3u
        MP817 N$5854 N$5897 N$5853 VDD p L=2u W=3u
        MP816 N$5853 N$4313 N$5852 VDD p L=2u W=3u
        MP820 OUT5 N$5855 VDD VDD p L=2u W=3u
        MN819 N$5855 N$5833 N$5857 GND n L=2u W=3u
        MN818 N$5855 N$5847 N$5856 GND n L=2u W=3u
        MN817 N$5858 N$5897 GND GND n L=2u W=3u
        MN816 N$5857 N$4313 N$5858 GND n L=2u W=3u
        MN815 N$5856 N$5833 GND GND n L=2u W=3u
        MP825 N$5863 N$4314 N$5862 VDD p L=2u W=3u
        MP824 N$5863 N$5849 N$5861 VDD p L=2u W=3u
        MP823 N$5862 N$5942 N$5861 VDD p L=2u W=3u
        MP822 N$5861 N$5942 VDD VDD p L=2u W=3u
        MP797 N$5831 N$4348 N$5830 VDD p L=2u W=3u
        MP796 N$5831 N$5817 N$5829 VDD p L=2u W=3u
        MP795 N$5830 N$5896 N$5829 VDD p L=2u W=3u
        MP794 N$5829 N$5896 VDD VDD p L=2u W=3u
        MP793 N$5829 N$4348 VDD VDD p L=2u W=3u
        MP798 N$5833 N$5831 VDD VDD p L=2u W=3u
        MN798 N$5831 N$4348 N$5835 GND n L=2u W=3u
        MN797 N$5834 N$5896 GND GND n L=2u W=3u
        MN796 N$5835 N$5896 GND GND n L=2u W=3u
        MP831 N$5870 N$5942 N$5869 VDD p L=2u W=3u
        MP830 N$5869 N$4314 N$5868 VDD p L=2u W=3u
        MP829 N$5868 N$5942 VDD VDD p L=2u W=3u
        MP828 N$5868 N$4314 VDD VDD p L=2u W=3u
        MP827 N$5868 N$5849 VDD VDD p L=2u W=3u
        MN831 N$5874 N$5942 GND GND n L=2u W=3u
        MN830 N$5873 N$4314 N$5874 GND n L=2u W=3u
        MN829 N$5872 N$5849 GND GND n L=2u W=3u
        MN828 N$5872 N$5942 GND GND n L=2u W=3u
        MN827 N$5872 N$4314 GND GND n L=2u W=3u
        MP833 N$5871 N$5863 N$5868 VDD p L=2u W=3u
        MP836 N$5877 N$5956 VDD VDD p L=2u W=3u
        MP835 N$5877 N$4315 VDD VDD p L=2u W=3u
        MN834 OUT6 N$5871 GND GND n L=2u W=3u
        MP834 OUT6 N$5871 VDD VDD p L=2u W=3u
        MN833 N$5871 N$5849 N$5873 GND n L=2u W=3u
        MN832 N$5871 N$5863 N$5872 GND n L=2u W=3u
        MN837 N$5879 N$5865 N$5882 GND n L=2u W=3u
        MN836 N$5882 N$4315 GND GND n L=2u W=3u
        MN805 N$5839 N$5817 N$5841 GND n L=2u W=3u
        MN804 N$5839 N$5831 N$5840 GND n L=2u W=3u
        MN809 N$5847 N$5833 N$5850 GND n L=2u W=3u
        MN808 N$5850 N$4313 GND GND n L=2u W=3u
        MN807 N$5849 N$5847 GND GND n L=2u W=3u
        MP811 N$5847 N$4313 N$5846 VDD p L=2u W=3u
        MP810 N$5847 N$5833 N$5845 VDD p L=2u W=3u
        MP809 N$5846 N$5897 N$5845 VDD p L=2u W=3u
        MP815 N$5852 N$5897 VDD VDD p L=2u W=3u
        MP814 N$5852 N$4313 VDD VDD p L=2u W=3u
        MP813 N$5852 N$5833 VDD VDD p L=2u W=3u
        MN842 N$5888 N$5956 GND GND n L=2u W=3u
        MN841 N$5888 N$4315 GND GND n L=2u W=3u
        MP847 N$5887 N$5879 N$5884 VDD p L=2u W=3u
        MP846 N$5887 N$5865 N$5886 VDD p L=2u W=3u
        MP845 N$5886 N$5956 N$5885 VDD p L=2u W=3u
        MP844 N$5885 N$4315 N$5884 VDD p L=2u W=3u
        MP848 OUT7 N$5887 VDD VDD p L=2u W=3u
        MN847 N$5887 N$5865 N$5889 GND n L=2u W=3u
        MN846 N$5887 N$5879 N$5888 GND n L=2u W=3u
        MN845 N$5890 N$5956 GND GND n L=2u W=3u
        MN844 N$5889 N$4315 N$5890 GND n L=2u W=3u
        MN843 N$5888 N$5865 GND GND n L=2u W=3u
        MP230 N$5969 CK N$5978 VDD p L=2u W=6u
        MN230 N$5978 N$5966 N$5969 GND n L=2u W=6u
        MP229 N$5967 N$5966 N$5969 VDD p L=2u W=6u
        MN229 N$5969 CK N$5967 GND n L=2u W=6u
        MN228 N$5967 N$5968 GND GND n L=2u W=6u
        MP228 N$5967 N$5968 VDD VDD p L=2u W=6u
        MP821 N$5861 N$4314 VDD VDD p L=2u W=3u
        MN820 OUT5 N$5855 GND GND n L=2u W=3u
        MP826 N$5865 N$5863 VDD VDD p L=2u W=3u
        MN826 N$5863 N$4314 N$5867 GND n L=2u W=3u
        MN825 N$5866 N$5942 GND GND n L=2u W=3u
        MN824 N$5867 N$5942 GND GND n L=2u W=3u
        MN823 N$5863 N$5849 N$5866 GND n L=2u W=3u
        MN822 N$5866 N$4314 GND GND n L=2u W=3u
        MN821 N$5865 N$5863 GND GND n L=2u W=3u
        MP832 N$5871 N$5849 N$5870 VDD p L=2u W=3u
        MN115 N$953 N$1579 GND GND n L=2u W=3u
        MN116 N$953 N$2908 GND GND n L=2u W=3u
        MP73 N$1032 N$6186 VDD VDD p L=2u W=6u
        MN72 N$1032 N$6186 N$1028 GND n L=2u W=6u
        MP72 N$1032 N$4990 VDD VDD p L=2u W=6u
        MN71 N$2907 N$1033 GND GND n L=2u W=6u
        MP138 N$1051 N$5204 VDD VDD p L=2u W=6u
        MP215 N$1068 N$5744 VDD VDD p L=2u W=6u
        MN214 N$1068 N$5744 N$1069 GND n L=2u W=6u
        MP214 N$1068 N$4989 VDD VDD p L=2u W=6u
        MN213 N$1607 N$1066 GND GND n L=2u W=6u
        MN96 N$933 N$1578 GND GND n L=2u W=3u
        MN95 N$2494 N$932 GND GND n L=2u W=3u
        MP99 N$932 N$1578 N$931 VDD p L=2u W=3u
        MP98 N$932 N$25 N$929 VDD p L=2u W=3u
        MP97 N$931 N$51 N$929 VDD p L=2u W=3u
        MP96 N$929 N$51 VDD VDD p L=2u W=3u
        MP95 N$929 N$1578 VDD VDD p L=2u W=3u
        MP120 N$952 N$41 N$951 VDD p L=2u W=3u
        MN122 N$956 N$952 GND GND n L=2u W=3u
        MN835 CARRY_OUT N$5879 GND GND n L=2u W=3u
        MP839 N$5879 N$4315 N$5878 VDD p L=2u W=3u
        MP838 N$5879 N$5865 N$5877 VDD p L=2u W=3u
        MP837 N$5878 N$5956 N$5877 VDD p L=2u W=3u
        MP843 N$5884 N$5956 VDD VDD p L=2u W=3u
        MP842 N$5884 N$4315 VDD VDD p L=2u W=3u
        MP841 N$5884 N$5865 VDD VDD p L=2u W=3u
        MP840 CARRY_OUT N$5879 VDD VDD p L=2u W=3u
        MN840 N$5879 N$4315 N$5883 GND n L=2u W=3u
        MN839 N$5882 N$5956 GND GND n L=2u W=3u
        MN838 N$5883 N$5956 GND GND n L=2u W=3u
        MP172 N$993 N$709 N$992 VDD p L=2u W=3u
        MP171 N$992 N$942 VDD VDD p L=2u W=3u
        MP170 N$992 N$709 VDD VDD p L=2u W=3u
        MP176 N$999 N$995 VDD VDD p L=2u W=3u
        MN175 N$995 N$2903 N$997 GND n L=2u W=3u
        MN174 N$995 N$988 N$996 GND n L=2u W=3u
        MN173 N$998 N$942 GND GND n L=2u W=3u
        MN172 N$997 N$709 N$998 GND n L=2u W=3u
        MN171 N$996 N$2903 GND GND n L=2u W=3u
        MP186 N$1007 N$2902 N$1006 VDD p L=2u W=3u
        MP185 N$1006 N$956 VDD VDD p L=2u W=3u
        MP174 N$995 N$2903 N$994 VDD p L=2u W=3u
        MN46 N$3666 N$3701 GND GND n L=2u W=3u
        MN45 N$3664 GND N$3665 GND n L=2u W=3u
        MN44 N$3665 N$3451 GND GND n L=2u W=3u
        MN43 N$3700 N$3664 GND GND n L=2u W=3u
        MP47 N$3664 N$3451 N$3663 VDD p L=2u W=3u
        MP46 N$3664 GND N$3662 VDD p L=2u W=3u
        MP45 N$3663 N$3701 N$3662 VDD p L=2u W=3u
        MP44 N$3662 N$3701 VDD VDD p L=2u W=3u
        MP43 N$3662 N$3451 VDD VDD p L=2u W=3u
        MN848 OUT7 N$5887 GND GND n L=2u W=3u
        MN227 N$5968 N$5965 GND GND n L=2u W=6u
        MP121 N$952 N$945 N$949 VDD p L=2u W=3u
        MP241 N$5979 N$5980 VDD VDD p L=2u W=6u
        MN240 N$5975 N$5979 GND GND n L=2u W=6u
        MP240 N$5975 N$5979 VDD VDD p L=2u W=6u
        MP239 N$5980 CK N$5975 VDD p L=2u W=6u
        MN239 N$5975 N$5983 N$5980 GND n L=2u W=6u
        MP238 N$5982 N$5983 N$5980 VDD p L=2u W=6u
        MN238 N$5980 CK N$5982 GND n L=2u W=6u
        MN237 N$5982 N$5981 GND GND n L=2u W=6u
        MP237 N$5982 N$5981 VDD VDD p L=2u W=6u
        MN236 N$5981 N$5984 GND GND n L=2u W=6u
        MP236 N$5981 N$5984 VDD VDD p L=2u W=6u
        MP235 N$5984 N$5983 N$5982 VDD p L=2u W=6u
        MN235 N$5982 CK N$5984 GND n L=2u W=6u
        MP234 N$5978 CK N$5984 VDD p L=2u W=6u
        MN234 N$5984 N$5983 N$5978 GND n L=2u W=6u
        MP233 N$5966 CK VDD VDD p L=2u W=5u
        MN233 N$5966 CK GND GND n L=2u W=5u
        MN232 N$5970 N$5969 GND GND n L=2u W=6u
        MP232 N$5970 N$5969 VDD VDD p L=2u W=6u
        MN231 N$5978 N$5970 GND GND n L=2u W=6u
        MP231 N$5978 N$5970 VDD VDD p L=2u W=6u
        MP122 N$956 N$952 VDD VDD p L=2u W=3u
        MN121 N$952 N$41 N$954 GND n L=2u W=3u
        MN120 N$952 N$945 N$953 GND n L=2u W=3u
        MN119 N$955 N$2908 GND GND n L=2u W=3u
        MN215 N$1069 N$4989 GND GND n L=2u W=6u
        MN16 N$26 N$2905 GND GND n L=2u W=3u
        MN15 N$25 N$24 GND GND n L=2u W=3u
        MP19 N$24 N$2905 N$23 VDD p L=2u W=3u
        MP18 N$24 GND N$20 VDD p L=2u W=3u
        MP227 N$5968 N$5965 VDD VDD p L=2u W=6u
        MP173 N$994 N$942 N$993 VDD p L=2u W=3u
        MP344 A0 N$5979 N$5920 VDD p L=2u W=5u
        MN343 N$5919 N$5979 GND GND n L=2u W=5u
        MP343 GND N$5958 N$5919 VDD p L=2u W=5u
        MN342 N$5919 N$5958 A1 GND n L=2u W=5u
        MP342 A1 N$5979 N$5919 VDD p L=2u W=5u
        MN341 N$5918 N$5979 GND GND n L=2u W=5u
        MP341 GND N$5958 N$5918 VDD p L=2u W=5u
        MN340 N$5918 N$5958 A2 GND n L=2u W=5u
        MN306 N$5983 CK GND GND n L=2u W=5u
        MP306 N$5983 CK VDD VDD p L=2u W=5u
        MN241 N$5979 N$5980 GND GND n L=2u W=6u
        MP614 N$5356 N$5358 VDD VDD p L=2u W=6u
        MN613 N$5357 N$5356 GND GND n L=2u W=6u
        MP613 N$5357 N$5356 VDD VDD p L=2u W=6u
        MP612 N$5358 CK N$5357 VDD p L=2u W=6u
        MN612 N$5357 N$5362 N$5358 GND n L=2u W=6u
        MP617 N$5355 N$5354 N$5352 VDD p L=2u W=6u
        MN617 N$5352 CK N$5355 GND n L=2u W=6u
        MP616 N$5353 CK N$5355 VDD p L=2u W=6u
        MN616 N$5355 N$5354 N$5353 GND n L=2u W=6u
        MN615 N$5362 CK GND GND n L=2u W=5u
        MN614 N$5356 N$5358 GND GND n L=2u W=6u
        MP615 N$5362 CK VDD VDD p L=2u W=5u
        MN621 N$5349 N$5354 N$5350 GND n L=2u W=6u
        MP620 N$5352 N$5354 N$5350 VDD p L=2u W=6u
        MN620 N$5350 CK N$5352 GND n L=2u W=6u
        MN619 N$5352 N$5351 GND GND n L=2u W=6u
        MP619 N$5352 N$5351 VDD VDD p L=2u W=6u
        MN618 N$5351 N$5355 GND GND n L=2u W=6u
        MP618 N$5351 N$5355 VDD VDD p L=2u W=6u
        MP670 N$5303 N$5310 N$5306 VDD p L=2u W=3u
        MP669 N$5303 N$5324 N$5304 VDD p L=2u W=3u
        MP681 N$5298 B2 VDD VDD p L=2u W=3u
        MN670 N$5299 N$5303 GND GND n L=2u W=3u
        MP671 N$5299 N$5303 VDD VDD p L=2u W=3u
        MN669 N$5303 N$5324 N$5301 GND n L=2u W=3u
        MN668 N$5303 N$5310 N$5302 GND n L=2u W=3u
        MN642 N$5333 N$5338 GND GND n L=2u W=5u
        MP642 GND N$5910 N$5333 VDD p L=2u W=5u
        MN466 N$5489 N$5492 N$5486 GND n L=2u W=3u
        MN465 N$5487 N$5491 GND GND n L=2u W=3u
        MN464 N$5486 N$5491 GND GND n L=2u W=3u
        MN463 N$5489 N$5505 N$5487 GND n L=2u W=3u
        MN462 N$5487 N$5492 GND GND n L=2u W=3u
        MP472 N$5482 N$5505 N$5483 VDD p L=2u W=3u
        MP471 N$5483 N$5491 N$5484 VDD p L=2u W=3u
        MP470 N$5484 N$5492 N$5485 VDD p L=2u W=3u
        MP469 N$5485 N$5491 VDD VDD p L=2u W=3u
        MP468 N$5485 N$5492 VDD VDD p L=2u W=3u
        MP467 N$5485 N$5505 VDD VDD p L=2u W=3u
        MN472 N$5482 N$5489 N$5481 GND n L=2u W=3u
        MP462 N$5493 N$5491 VDD VDD p L=2u W=3u
        MN470 N$5480 N$5492 N$5479 GND n L=2u W=3u
        MN469 N$5481 N$5505 GND GND n L=2u W=3u
        MN468 N$5481 N$5491 GND GND n L=2u W=3u
        MN467 N$5481 N$5492 GND GND n L=2u W=3u
        MP473 N$5482 N$5489 N$5485 VDD p L=2u W=3u
        MP477 N$5476 N$5474 VDD VDD p L=2u W=3u
        MP476 N$5476 N$5475 VDD VDD p L=2u W=3u
        MN412 N$5937 N$5932 N$5928 GND n L=2u W=5u
        MP412 N$5928 N$5349 N$5937 VDD p L=2u W=5u
        MN411 N$5936 N$5349 N$5929 GND n L=2u W=5u
        MP411 N$5929 N$5932 N$5936 VDD p L=2u W=5u
        MN410 N$5936 N$5932 N$5927 GND n L=2u W=5u
        MP410 N$5927 N$5349 N$5936 VDD p L=2u W=5u
        MN409 N$5935 N$5349 N$5928 GND n L=2u W=5u
        MP409 N$5928 N$5932 N$5935 VDD p L=2u W=5u
        MP466 N$5488 N$5489 VDD VDD p L=2u W=3u
        MP625 N$5345 CK N$5347 VDD p L=2u W=6u
        MN625 N$5347 N$5346 N$5345 GND n L=2u W=6u
        MN624 N$5354 CK GND GND n L=2u W=5u
        MP630 N$5342 CK N$5341 VDD p L=2u W=6u
        MN630 N$5341 N$5346 N$5342 GND n L=2u W=6u
        MP629 N$5344 N$5346 N$5342 VDD p L=2u W=6u
        MN629 N$5342 CK N$5344 GND n L=2u W=6u
        MN628 N$5344 N$5343 GND GND n L=2u W=6u
        MP628 N$5344 N$5343 VDD VDD p L=2u W=6u
        MN627 N$5343 N$5347 GND GND n L=2u W=6u
        MN633 N$5346 CK GND GND n L=2u W=5u
        MN626 N$5344 CK N$5347 GND n L=2u W=6u
        MP633 N$5346 CK VDD VDD p L=2u W=5u
        MN632 N$5340 N$5342 GND GND n L=2u W=6u
        MP632 N$5340 N$5342 VDD VDD p L=2u W=6u
        MN631 N$5341 N$5340 GND GND n L=2u W=6u
        MP631 N$5341 N$5340 VDD VDD p L=2u W=6u
        MN636 N$5338 N$5910 GND GND n L=2u W=5u
        MP636 N$5338 N$5910 VDD VDD p L=2u W=5u
        MN635 N$5337 N$5338 GND GND n L=2u W=5u
        MP635 GND N$5910 N$5337 VDD p L=2u W=5u
        MN634 N$5337 N$5910 N$5420 GND n L=2u W=5u
        MN360 N$5928 N$5357 N$5919 GND n L=2u W=5u
        MP360 N$5919 N$5923 N$5928 VDD p L=2u W=5u
        MN359 N$5928 N$5923 N$5918 GND n L=2u W=5u
        MP359 N$5918 N$5357 N$5928 VDD p L=2u W=5u
        MN358 N$5927 N$5357 N$5918 GND n L=2u W=5u
        MP358 N$5918 N$5923 N$5927 VDD p L=2u W=5u
        MN357 N$5927 N$5923 N$5917 GND n L=2u W=5u
        MP357 N$5917 N$5357 N$5927 VDD p L=2u W=5u
        MN424 N$5897 N$5341 N$5937 GND n L=2u W=5u
        MP424 N$5937 N$5941 N$5897 VDD p L=2u W=5u
        MN423 N$5897 N$5941 N$5934 GND n L=2u W=5u



*.ends mynand3

* Auxiliary circuit for power analysis
Cp Pav 0 100p
Rp Pav 0 100k
Fp 0 Pav Vtstp 0.003125
*Output load capacitance if you have any

*Cload1 out GND 200fF
.MODEL n NMOS LEVEL = 3
+ TOX = 200E-10 NSUB = 1E17 GAMMA = 0.5
+ PHI = 0.7 VTO = 0.8 DELTA = 3.0
+ UO = 650 ETA = 3.0E-6 THETA = 0.1
+ KP = 120E-6 VMAX = 1E5 KAPPA = 0.3
+ RSH = 0 NFS = 1E12 TPG = 1
+ XJ = 500E-9 LD = 100E-9
+ CGDO = 200E-12 CGSO = 200E-12 CGBO = 1E-10
+ CJ = 400E-6 PB = 1 MJ = 0.5
+ CJSW = 300E-12 MJSW = 0.5

.MODEL p PMOS LEVEL = 3
+ TOX = 200E-10 NSUB = 1E17 GAMMA = 0.6
+ PHI = 0.7 VTO = -0.9 DELTA = 0.1
+ UO = 250 ETA = 0 THETA = 0.1
+ KP = 40E-6 VMAX = 5E4 KAPPA = 1
+ RSH = 0 NFS = 1E12 TPG = -1
+ XJ = 500E-9 LD = 100E-9
+ CGDO = 200E-12 CGSO = 200E-12 CGBO = 1E-10
+ CJ = 400E-6 PB = 1 MJ = 0.5
+ CJSW = 300E-12 MJSW = 0.5

*Define power rails
Vddt top 0 5
Vtstp top Vdd 0
Vss GND 0 0

* Define input voltages of A and B

Vck CK 0 PWL(0 5 20N 5 20.1N 0 40N 0 40.1N 5 60N 5 60.1N 0 80N 0 80.1N 5 100N 5 
+ 100.1N 0 120N 0 120.1N 5 140N 5 140.1N 0 160N 0 160.1N 5 180N 5 180.1N 0 200N 0
+ 200.1N 5 220N 5 220.1N 0 240N 0 240.1N 5 260N 5 260.1N 0 280N 0 280.1N 5 300N 5 
+ 300.1N 0 320N 0 320.1N 5 340N 5 340.1N 0 360N 0 360.1N 5 380N 5 380.1N 0 400N 0 
+ 400.1N 0 420N 0 420.1N 5 440N 5 440.1N 0 460N 0 460.1N 5 480N 5 480.1N 0 500N 0)
Va5 A5 0 PWL(0 5 20N 5 20.1N 5 40N 5 40.1N 0 60N 0 60.1N 0 80N 0 80.1N 0 100N 0 
+ 100.1N 0 120N 0 120.1N 0 140N 0 140.1N 0 160N 0 160.1N 0 180N 0 180.1N 0 200N 0
+ 200.1N 0 220N 0 220.1N 0 240N 0 240.1N 0 260N 0 260.1N 0 280N 0 280.1N 0 300N 0 
+ 300.1N 0 320N 0 320.1N 0 340N 0 340.1N 0 360N 0 360.1N 0 380N 0 380.1N 0 400N 0 
+ 400.1N 0 420N 0 420.1N 0 440N 0 440.1N 0 460N 0 460.1N 0 480N 0 480.1N 0 500N 0)
Va0 A0 0 PWL(0 5 20N 5 20.1N 5 40N 5 40.1N 5 60N 5 60.1N 5 80N 5 80.1N 5 100N 5 
+ 100.1N 5 120N 5 120.1N 5 140N 5 140.1N 5 160N 5 160.1N 5 180N 5 180.1N 5 200N 5
+ 200.1N 5 220N 5 220.1N 5 240N 5 240.1N 5 260N 5 260.1N 5 280N 5 280.1N 5 300N 5 
+ 300.1N 5 320N 5 320.1N 5 340N 5 340.1N 5 360N 5 360.1N 5 380N 5 380.1N 5 400N 5 
+ 400.1N 5 420N 5 420.1N 5 440N 5 440.1N 5 460N 5 460.1N 5 480N 5 480.1N 5 500N 5)
Va2 A2 0 PWL(0 0 20N 0 20.1N 0 40N 0 40.1N 0 60N 0 60.1N 0 80N 0 80.1N 0 100N 0 
+ 100.1N 0 120N 0 120.1N 0 140N 0 140.1N 0 160N 0 160.1N 0 180N 0 180.1N 0 200N 0
+ 200.1N 0 220N 0 220.1N 0 240N 0 240.1N 0 260N 0 260.1N 0 280N 0 280.1N 0 300N 0 
+ 300.1N 0 320N 0 320.1N 0 340N 0 340.1N 0 360N 0 360.1N 0 380N 0 380.1N 0 400N 0 
+ 400.1N 0 420N 0 420.1N 0 440N 0 440.1N 0 460N 0 460.1N 0 480N 0 480.1N 0 500N 0)
Va1 A1 0 PWL(0 5 20N 5 20.1N 5 40N 5 40.1N 5 60N 5 60.1N 5 80N 5 80.1N 5 100N 5 
+ 100.1N 5 120N 5 120.1N 5 140N 5 140.1N 5 160N 5 160.1N 5 180N 5 180.1N 5 200N 5
+ 200.1N 5 220N 5 220.1N 5 240N 5 240.1N 5 260N 5 260.1N 5 280N 5 280.1N 5 300N 5 
+ 300.1N 5 320N 5 320.1N 5 340N 5 340.1N 5 360N 5 360.1N 5 380N 5 380.1N 5 400N 5 
+ 400.1N 5 420N 5 420.1N 5 440N 5 440.1N 5 460N 5 460.1N 5 480N 5 480.1N 5 500N 5)
Va3 A3 0 PWL(0 0 20N 0 20.1N 0 40N 0 40.1N 0 60N 0 60.1N 0 80N 0 80.1N 0 100N 0 
+ 100.1N 0 120N 0 120.1N 0 140N 0 140.1N 0 160N 0 160.1N 0 180N 0 180.1N 0 200N 0
+ 200.1N 0 220N 0 220.1N 0 240N 0 240.1N 0 260N 0 260.1N 0 280N 0 280.1N 0 300N 0 
+ 300.1N 0 320N 0 320.1N 0 340N 0 340.1N 0 360N 0 360.1N 0 380N 0 380.1N 0 400N 0 
+ 400.1N 0 420N 0 420.1N 0 440N 0 440.1N 0 460N 0 460.1N 0 480N 0 480.1N 0 500N 0)
Vrst RST 0 PWL(0 5 20N 5 20.1N 5 40N 5 40.1N 0 60N 0 60.1N 0 80N 0 80.1N 0 100N 0 
+ 100.1N 0 120N 0 120.1N 0 140N 0 140.1N 0 160N 0 160.1N 0 180N 0 180.1N 0 200N 0
+ 200.1N 0 220N 0 220.1N 0 240N 0 240.1N 0 260N 0 260.1N 0 280N 0 280.1N 0 300N 0 
+ 300.1N 0 320N 0 320.1N 0 340N 0 340.1N 0 360N 0 360.1N 0 380N 0 380.1N 0 400N 0 
+ 400.1N 0 420N 0 420.1N 0 440N 0 440.1N 0 460N 0 460.1N 0 480N 0 480.1N 0 500N 0)
Vb0 B0 0 PWL(0 5 20N 5 20.1N 5 40N 5 40.1N 5 60N 5 60.1N 5 80N 5 80.1N 5 100N 5 
+ 100.1N 5 120N 5 120.1N 5 140N 5 140.1N 5 160N 5 160.1N 5 180N 5 180.1N 5 200N 5
+ 200.1N 5 220N 5 220.1N 5 240N 5 240.1N 5 260N 5 260.1N 5 280N 5 280.1N 5 300N 5 
+ 300.1N 5 320N 5 320.1N 5 340N 5 340.1N 5 360N 5 360.1N 5 380N 5 380.1N 5 400N 5 
+ 400.1N 5 420N 5 420.1N 5 440N 5 440.1N 5 460N 5 460.1N 5 480N 5 480.1N 5 500N 5)
Vb1 B1 0 PWL(0 0 20N 0 20.1N 0 40N 0 40.1N 0 60N 0 60.1N 0 80N 0 80.1N 0 100N 0 
+ 100.1N 0 120N 0 120.1N 0 140N 0 140.1N 0 160N 0 160.1N 0 180N 0 180.1N 0 200N 0
+ 200.1N 0 220N 0 220.1N 0 240N 0 240.1N 0 260N 0 260.1N 0 280N 0 280.1N 0 300N 0 
+ 300.1N 0 320N 0 320.1N 0 340N 0 340.1N 0 360N 0 360.1N 0 380N 0 380.1N 0 400N 0 
+ 400.1N 0 420N 0 420.1N 0 440N 0 440.1N 0 460N 0 460.1N 0 480N 0 480.1N 0 500N 0)
Vb2 B2 0 PWL(0 5 20N 5 20.1N 5 40N 5 40.1N 5 60N 5 60.1N 5 80N 5 80.1N 5 100N 5 
+ 100.1N 5 120N 5 120.1N 5 140N 5 140.1N 5 160N 5 160.1N 5 180N 5 180.1N 5 200N 5
+ 200.1N 5 220N 5 220.1N 5 240N 5 240.1N 5 260N 5 260.1N 5 280N 5 280.1N 5 300N 5 
+ 300.1N 5 320N 5 320.1N 5 340N 5 340.1N 5 360N 5 360.1N 5 380N 5 380.1N 5 400N 5 
+ 400.1N 5 420N 5 420.1N 5 440N 5 440.1N 5 460N 5 460.1N 5 480N 5 480.1N 5 500N 5)
Vb3 B3 0 PWL(0 0 20N 0 20.1N 0 40N 0 40.1N 0 60N 0 60.1N 0 80N 0 80.1N 0 100N 0 
+ 100.1N 0 120N 0 120.1N 0 140N 0 140.1N 0 160N 0 160.1N 0 180N 0 180.1N 0 200N 0
+ 200.1N 0 220N 0 220.1N 0 240N 0 240.1N 0 260N 0 260.1N 0 280N 0 280.1N 0 300N 0 
+ 300.1N 0 320N 0 320.1N 0 340N 0 340.1N 0 360N 0 360.1N 0 380N 0 380.1N 0 400N 0 
+ 400.1N 0 420N 0 420.1N 0 440N 0 440.1N 0 460N 0 460.1N 0 480N 0 480.1N 0 500N 0)
Vc C 0 PWL(0 0 20N 0 20.1N 0 40N 0 40.1N 0 60N 0 60.1N 0 80N 0 80.1N 0 100N 0 
+ 100.1N 0 120N 0 120.1N 0 140N 0 140.1N 0 160N 0 160.1N 0 180N 0 180.1N 0 200N 0
+ 200.1N 0 220N 0 220.1N 0 240N 0 240.1N 0 260N 0 260.1N 0 280N 0 280.1N 0 300N 0 
+ 300.1N 0 320N 0 320.1N 0 340N 0 340.1N 0 360N 0 360.1N 0 380N 0 380.1N 0 400N 0 
+ 400.1N 0 420N 0 420.1N 0 440N 0 440.1N 0 460N 0 460.1N 0 480N 0 480.1N 0 500N 0)



*Define transient simulation and probe voltage/current signals
.TRAN 20N 500N
.PROBE V(*) I(*)
.end
