




*.subckt mynand3 A B GND Out Vdd



* MAIN CELL: Component pathname : /home/mentor/jack/jaggu
*
        MP280 N$4357 N$4360 N$4356 VDD p L=2u W=6u
        MP281 N$4359 N$4357 VDD VDD p L=2u W=6u
        MN281 N$4359 N$4357 GND GND n L=2u W=6u
        MP282 N$4356 N$4359 VDD VDD p L=2u W=6u
        MN282 N$4356 N$4359 GND GND n L=2u W=6u
        MN283 N$4355 CLK N$4356 GND n L=2u W=6u
        MP283 N$4356 N$4360 N$4355 VDD p L=2u W=6u
        MN284 P5 N$4360 N$4355 GND n L=2u W=6u
        MP284 N$4355 CLK P5 VDD p L=2u W=6u
        MP285 P5 N$4358 VDD VDD p L=2u W=6u
        MN285 P5 N$4358 GND GND n L=2u W=6u
        MP286 N$4358 N$4355 VDD VDD p L=2u W=6u
        MN144 N$1058 B2 GND GND n L=2u W=6u
        MN212 N$1067 B2 GND GND n L=2u W=6u
        MP144 N$1057 A2 VDD VDD p L=2u W=6u
        MN209 N$1065 B0 GND GND n L=2u W=6u
        MP209 N$1064 A3 VDD VDD p L=2u W=6u
        MN208 N$1064 A3 N$1065 GND n L=2u W=6u
        MP208 N$1064 B0 VDD VDD p L=2u W=6u
        MN207 N$2902 N$1077 GND GND n L=2u W=6u
        MP167 N$988 N$709 N$987 VDD p L=2u W=3u
        MP28 N$1601 N$31 VDD VDD p L=2u W=3u
        MN34 N$40 N$2904 N$43 GND n L=2u W=3u
        MN33 N$42 N$2906 GND GND n L=2u W=3u
        MN32 N$43 N$2906 GND GND n L=2u W=3u
        MN31 N$40 C1 N$42 GND n L=2u W=3u
        MN30 N$42 N$2904 GND GND n L=2u W=3u
        MN29 N$41 N$40 GND GND n L=2u W=3u
        MP33 N$40 N$2904 N$39 VDD p L=2u W=3u
        MP39 N$46 N$2906 N$45 VDD p L=2u W=3u
        MP38 N$45 N$2904 N$44 VDD p L=2u W=3u
        MP37 N$44 N$2906 VDD VDD p L=2u W=3u
        MP132 N$3681 N$2491 N$3680 VDD p L=2u W=3u
        MP131 N$3680 N$3446 VDD VDD p L=2u W=3u
        MP130 N$3680 N$2491 VDD VDD p L=2u W=3u
        MP129 N$3680 N$3700 VDD VDD p L=2u W=3u
        MP128 N$3460 N$3677 VDD VDD p L=2u W=3u
        MN128 N$3677 N$2491 N$3679 GND n L=2u W=3u
        MN127 N$3678 N$3446 GND GND n L=2u W=3u
        MN126 N$3679 N$3446 GND GND n L=2u W=3u
        MN125 N$3677 N$3700 N$3678 GND n L=2u W=3u
        MN124 N$3678 N$2491 GND GND n L=2u W=3u
        MN123 N$3460 N$3677 GND GND n L=2u W=3u
        MP126 N$3677 N$3700 N$3675 VDD p L=2u W=3u
        MN3 N$6 C1 N$10 GND n L=2u W=3u
        MN2 N$10 N$4109 GND GND n L=2u W=3u
        MN1 N$9 N$6 GND GND n L=2u W=3u
        MP125 N$3676 N$3446 N$3675 VDD p L=2u W=3u
        MP124 N$3675 N$3446 VDD VDD p L=2u W=3u
        MP123 N$3675 N$2491 VDD VDD p L=2u W=3u
        MN135 N$3683 N$3700 N$3685 GND n L=2u W=3u
        MN56 N$4320 N$3670 GND GND n L=2u W=3u
        MP56 N$4320 N$3670 VDD VDD p L=2u W=3u
        MP127 N$3677 N$2491 N$3676 VDD p L=2u W=3u
        MP117 N$949 N$2908 VDD VDD p L=2u W=3u
        MP118 N$950 N$1579 N$949 VDD p L=2u W=3u
        MN73 N$1028 B0 GND GND n L=2u W=6u
        MN13 N$15 C1 N$17 GND n L=2u W=3u
        MN12 N$15 N$6 N$16 GND n L=2u W=3u
        MN11 N$18 N$2907 GND GND n L=2u W=3u
        MP116 N$949 N$1579 VDD VDD p L=2u W=3u
        MP5 N$6 N$4109 N$5 VDD p L=2u W=3u
        MP4 N$6 C1 N$2 VDD p L=2u W=3u
        MP157 N$3693 N$3456 VDD VDD p L=2u W=3u
        MP244 N$4331 N$4334 N$4330 VDD p L=2u W=6u
        MN244 N$4330 CLK N$4331 GND n L=2u W=6u
        MP243 N$2020 CLK N$4331 VDD p L=2u W=6u
        MN243 N$4331 N$4334 N$2020 GND n L=2u W=6u
        MN242 N$4328 CLK GND GND n L=2u W=5u
        MP242 N$4328 CLK VDD VDD p L=2u W=5u
        MN224 N$4326 N$4323 GND GND n L=2u W=6u
        MP224 N$4326 N$4323 VDD VDD p L=2u W=6u
        MN223 P0 N$4326 GND GND n L=2u W=6u
        MP223 P0 N$4326 VDD VDD p L=2u W=6u
        MP222 N$4323 CLK P0 VDD p L=2u W=6u
        MN222 P0 N$4328 N$4323 GND n L=2u W=6u
        MN300 N$4368 N$4371 GND GND n L=2u W=6u
        MP300 N$4368 N$4371 VDD VDD p L=2u W=6u
        MN299 N$4371 N$4369 GND GND n L=2u W=6u
        MP299 N$4371 N$4369 VDD VDD p L=2u W=6u
        MP298 N$4369 N$4372 N$4368 VDD p L=2u W=6u
        MN298 N$4368 CLK N$4369 GND n L=2u W=6u
        MP297 N$3690 CLK N$4369 VDD p L=2u W=6u
        MN297 N$4369 N$4372 N$3690 GND n L=2u W=6u
        MN296 N$4366 CLK GND GND n L=2u W=5u
        MP296 N$4366 CLK VDD VDD p L=2u W=5u
        MN301 N$4367 CLK N$4368 GND n L=2u W=6u
        MN134 N$3683 N$3677 N$3684 GND n L=2u W=3u
        MN133 N$3686 N$3446 GND GND n L=2u W=3u
        MN132 N$3685 N$2491 N$3686 GND n L=2u W=3u
        MN131 N$3684 N$3700 GND GND n L=2u W=3u
        MN130 N$3684 N$3446 GND GND n L=2u W=3u
        MN129 N$3684 N$2491 GND GND n L=2u W=3u
        MP135 N$3683 N$3677 N$3680 VDD p L=2u W=3u
        MP134 N$3683 N$3700 N$3682 VDD p L=2u W=3u
        MP133 N$3682 N$3446 N$3681 VDD p L=2u W=3u
        MN107 N$938 N$25 N$940 GND n L=2u W=3u
        MN106 N$938 N$932 N$939 GND n L=2u W=3u
        MN105 N$941 N$51 GND GND n L=2u W=3u
        MP141 N$1055 A2 VDD VDD p L=2u W=6u
        MN140 N$1055 A2 N$1056 GND n L=2u W=6u
        MP140 N$1055 B0 VDD VDD p L=2u W=6u
        MN139 N$1578 N$1051 GND GND n L=2u W=6u
        MP86 N$2903 N$916 VDD VDD p L=2u W=3u
        MN86 N$916 N$707 N$920 GND n L=2u W=3u
        MP87 N$921 N$9 VDD VDD p L=2u W=3u
        MP88 N$921 N$707 VDD VDD p L=2u W=3u
        MP89 N$921 N$1601 VDD VDD p L=2u W=3u
        MP90 N$922 N$707 N$921 VDD p L=2u W=3u
        MN195 N$1018 N$1584 GND GND n L=2u W=3u
        MN194 N$1019 N$1584 GND GND n L=2u W=3u
        MN197 N$1024 N$1607 GND GND n L=2u W=3u
        MP203 N$1023 N$1016 N$1020 VDD p L=2u W=3u
        MP202 N$1023 N$946 N$1022 VDD p L=2u W=3u
        MP201 N$1022 N$1584 N$1021 VDD p L=2u W=3u
        MP200 N$1021 N$1607 N$1020 VDD p L=2u W=3u
        MP199 N$1020 N$1584 VDD VDD p L=2u W=3u
        MN203 N$1023 N$946 N$1025 GND n L=2u W=3u
        MN202 N$1023 N$1016 N$1024 GND n L=2u W=3u
        MN201 N$1026 N$1584 GND GND n L=2u W=3u
        MN200 N$1025 N$1607 N$1026 GND n L=2u W=3u
        MN199 N$1024 N$946 GND GND n L=2u W=3u
        MN198 N$1024 N$1584 GND GND n L=2u W=3u
        MN103 N$939 N$25 GND GND n L=2u W=3u
        MN102 N$939 N$51 GND GND n L=2u W=3u
        MN101 N$939 N$1578 GND GND n L=2u W=3u
        MN196 N$1016 N$1607 N$1019 GND n L=2u W=3u
        MN206 N$1062 B1 GND GND n L=2u W=6u
        MP174 N$995 N$2903 N$994 VDD p L=2u W=3u
        MP173 N$994 N$942 N$993 VDD p L=2u W=3u
        MP172 N$993 N$709 N$992 VDD p L=2u W=3u
        MP171 N$992 N$942 VDD VDD p L=2u W=3u
        MP170 N$992 N$709 VDD VDD p L=2u W=3u
        MP176 N$999 N$995 VDD VDD p L=2u W=3u
        MN175 N$995 N$2903 N$997 GND n L=2u W=3u
        MN174 N$995 N$988 N$996 GND n L=2u W=3u
        MN173 N$998 N$942 GND GND n L=2u W=3u
        MN172 N$997 N$709 N$998 GND n L=2u W=3u
        MN171 N$996 N$2903 GND GND n L=2u W=3u
        MP186 N$1007 N$2902 N$1006 VDD p L=2u W=3u
        MP185 N$1006 N$956 VDD VDD p L=2u W=3u
        MN46 N$3666 N$3701 GND GND n L=2u W=3u
        MN45 N$3664 C1 N$3665 GND n L=2u W=3u
        MN44 N$3665 N$3451 GND GND n L=2u W=3u
        MN43 N$3700 N$3664 GND GND n L=2u W=3u
        MP47 N$3664 N$3451 N$3663 VDD p L=2u W=3u
        MP46 N$3664 C1 N$3662 VDD p L=2u W=3u
        MP45 N$3663 N$3701 N$3662 VDD p L=2u W=3u
        MP44 N$3662 N$3701 VDD VDD p L=2u W=3u
        MP43 N$3662 N$3451 VDD VDD p L=2u W=3u
        MP188 N$1009 N$2494 N$1008 VDD p L=2u W=3u
        MP187 N$1008 N$956 N$1007 VDD p L=2u W=3u
        MN183 N$1010 N$2902 GND GND n L=2u W=3u
        MP189 N$1009 N$1002 N$1006 VDD p L=2u W=3u
        MP82 N$914 N$1601 VDD VDD p L=2u W=3u
        MP81 N$914 N$707 VDD VDD p L=2u W=3u
        MN89 N$925 N$9 GND GND n L=2u W=3u
        MN108 N$942 N$938 GND GND n L=2u W=3u
        MP108 N$942 N$938 VDD VDD p L=2u W=3u
        MN90 N$926 N$707 N$927 GND n L=2u W=3u
        MP104 N$936 N$1578 N$935 VDD p L=2u W=3u
        MP32 N$40 C1 N$36 VDD p L=2u W=3u
        MP31 N$39 N$2906 N$36 VDD p L=2u W=3u
        MP165 N$987 N$942 N$986 VDD p L=2u W=3u
        MP164 N$986 N$942 VDD VDD p L=2u W=3u
        MP163 N$986 N$709 VDD VDD p L=2u W=3u
        MN39 N$50 N$2906 GND GND n L=2u W=3u
        MP207 N$2902 N$1077 VDD VDD p L=2u W=6u
        MP8 N$12 N$4109 VDD VDD p L=2u W=3u
        MP11 N$14 N$2907 N$13 VDD p L=2u W=3u
        MP7 N$12 C1 VDD VDD p L=2u W=3u
        MN8 N$16 N$2907 GND GND n L=2u W=3u
        MN181 N$1004 N$956 GND GND n L=2u W=3u
        MN180 N$1005 N$956 GND GND n L=2u W=3u
        MN179 N$1002 N$2494 N$1004 GND n L=2u W=3u
        MN178 N$1004 N$2902 GND GND n L=2u W=3u
        MN177 N$3446 N$1002 GND GND n L=2u W=3u
        MP166 N$988 N$2903 N$986 VDD p L=2u W=3u
        MN191 N$1017 N$1016 GND GND n L=2u W=3u
        MP181 N$1002 N$2902 N$1001 VDD p L=2u W=3u
        MP180 N$1002 N$2494 N$1000 VDD p L=2u W=3u
        MP179 N$1001 N$956 N$1000 VDD p L=2u W=3u
        MP178 N$1000 N$956 VDD VDD p L=2u W=3u
        MP177 N$1000 N$2902 VDD VDD p L=2u W=3u
        MN163 N$3701 N$988 GND GND n L=2u W=3u
        MN164 N$990 N$709 GND GND n L=2u W=3u
        MN167 N$990 N$942 GND GND n L=2u W=3u
        MN166 N$991 N$942 GND GND n L=2u W=3u
        MN170 N$996 N$942 GND GND n L=2u W=3u
        MN169 N$996 N$709 GND GND n L=2u W=3u
        MP175 N$995 N$988 N$992 VDD p L=2u W=3u
        MN210 N$709 N$1064 GND GND n L=2u W=6u
        MP210 N$709 N$1064 VDD VDD p L=2u W=6u
        MN28 N$1601 N$31 GND GND n L=2u W=3u
        MP29 N$36 N$2904 VDD VDD p L=2u W=3u
        MP30 N$36 N$2906 VDD VDD p L=2u W=3u
        MP103 N$935 N$51 VDD VDD p L=2u W=3u
        MP102 N$935 N$1578 VDD VDD p L=2u W=3u
        MP101 N$935 N$25 VDD VDD p L=2u W=3u
        MP100 N$2494 N$932 VDD VDD p L=2u W=3u
        MN100 N$932 N$1578 N$934 GND n L=2u W=3u
        MN99 N$933 N$51 GND GND n L=2u W=3u
        MN98 N$934 N$51 GND GND n L=2u W=3u
        MN97 N$932 N$25 N$933 GND n L=2u W=3u
        MP184 N$1006 N$2902 VDD VDD p L=2u W=3u
        MP183 N$1006 N$2494 VDD VDD p L=2u W=3u
        MP182 N$3446 N$1002 VDD VDD p L=2u W=3u
        MN204 N$2491 N$1023 GND GND n L=2u W=3u
        MP204 N$2491 N$1023 VDD VDD p L=2u W=3u
        MN182 N$1002 N$2902 N$1005 GND n L=2u W=3u
        MN85 N$919 N$1601 GND GND n L=2u W=3u
        MN84 N$920 N$1601 GND GND n L=2u W=3u
        MN83 N$916 N$9 N$919 GND n L=2u W=3u
        MN82 N$919 N$707 GND GND n L=2u W=3u
        MN81 N$2903 N$916 GND GND n L=2u W=3u
        MP85 N$916 N$707 N$915 VDD p L=2u W=3u
        MP84 N$916 N$9 N$914 VDD p L=2u W=3u
        MP83 N$915 N$1601 N$914 VDD p L=2u W=3u
        MN118 N$954 N$1579 N$955 GND n L=2u W=3u
        MN117 N$953 N$41 GND GND n L=2u W=3u
        MN93 N$924 N$9 N$926 GND n L=2u W=3u
        MN92 N$924 N$916 N$925 GND n L=2u W=3u
        MN91 N$927 N$1601 GND GND n L=2u W=3u
        MP17 N$23 N$2017 N$20 VDD p L=2u W=3u
        MP16 N$20 N$2017 VDD VDD p L=2u W=3u
        MP15 N$20 N$2905 VDD VDD p L=2u W=3u
        MP21 N$28 C1 VDD VDD p L=2u W=3u
        MP20 N$25 N$24 VDD VDD p L=2u W=3u
        MN20 N$24 N$2905 N$27 GND n L=2u W=3u
        MN19 N$26 N$2017 GND GND n L=2u W=3u
        MN18 N$27 N$2017 GND GND n L=2u W=3u
        MN17 N$24 C1 N$26 GND n L=2u W=3u
        MP27 N$31 N$24 N$28 VDD p L=2u W=3u
        MP26 N$31 C1 N$30 VDD p L=2u W=3u
        MP25 N$30 N$2017 N$29 VDD p L=2u W=3u
        MP24 N$29 N$2905 N$28 VDD p L=2u W=3u
        MN7 N$16 N$4109 GND GND n L=2u W=3u
        MP13 N$15 N$6 N$12 VDD p L=2u W=3u
        MP12 N$15 C1 N$14 VDD p L=2u W=3u
        MN9 N$16 C1 GND GND n L=2u W=3u
        MN10 N$17 N$4109 N$18 GND n L=2u W=3u
        MP10 N$13 N$4109 N$12 VDD p L=2u W=3u
        MP9 N$12 N$2907 VDD VDD p L=2u W=3u
        MN41 N$47 C1 N$49 GND n L=2u W=3u
        MN40 N$47 N$40 N$48 GND n L=2u W=3u
        MP42 N$51 N$47 VDD VDD p L=2u W=3u
        MN42 N$51 N$47 GND GND n L=2u W=3u
        MP169 N$992 N$2903 VDD VDD p L=2u W=3u
        MP168 N$3701 N$988 VDD VDD p L=2u W=3u
        MN168 N$988 N$709 N$991 GND n L=2u W=3u
        MP40 N$47 C1 N$46 VDD p L=2u W=3u
        MN21 N$32 N$2905 GND GND n L=2u W=3u
        MP212 N$1066 A3 VDD VDD p L=2u W=6u
        MN211 N$1066 A3 N$1067 GND n L=2u W=6u
        MP211 N$1066 B2 VDD VDD p L=2u W=6u
        MP120 N$952 N$41 N$951 VDD p L=2u W=3u
        MP121 N$952 N$945 N$949 VDD p L=2u W=3u
        MN115 N$953 N$1579 GND GND n L=2u W=3u
        MN116 N$953 N$2908 GND GND n L=2u W=3u
        MP73 N$1032 A0 VDD VDD p L=2u W=6u
        MN72 N$1032 A0 N$1028 GND n L=2u W=6u
        MP72 N$1032 B0 VDD VDD p L=2u W=6u
        MN71 N$2907 N$1033 GND GND n L=2u W=6u
        MP138 N$1051 A2 VDD VDD p L=2u W=6u
        MP215 N$1068 A3 VDD VDD p L=2u W=6u
        MN214 N$1068 A3 N$1069 GND n L=2u W=6u
        MP214 N$1068 B3 VDD VDD p L=2u W=6u
        MN213 N$1607 N$1066 GND GND n L=2u W=6u
        MN96 N$933 N$1578 GND GND n L=2u W=3u
        MN95 N$2494 N$932 GND GND n L=2u W=3u
        MP99 N$932 N$1578 N$931 VDD p L=2u W=3u
        MP98 N$932 N$25 N$929 VDD p L=2u W=3u
        MP97 N$931 N$51 N$929 VDD p L=2u W=3u
        MP96 N$929 N$51 VDD VDD p L=2u W=3u
        MP95 N$929 N$1578 VDD VDD p L=2u W=3u
        MN122 N$956 N$952 GND GND n L=2u W=3u
        MP122 N$956 N$952 VDD VDD p L=2u W=3u
        MN121 N$952 N$41 N$954 GND n L=2u W=3u
        MN120 N$952 N$945 N$953 GND n L=2u W=3u
        MN119 N$955 N$2908 GND GND n L=2u W=3u
        MN215 N$1069 B3 GND GND n L=2u W=6u
        MN16 N$26 N$2905 GND GND n L=2u W=3u
        MN15 N$25 N$24 GND GND n L=2u W=3u
        MP19 N$24 N$2905 N$23 VDD p L=2u W=3u
        MP18 N$24 C1 N$20 VDD p L=2u W=3u
        MP66 N$1049 B3 VDD VDD p L=2u W=6u
        MN65 N$2904 N$1046 GND GND n L=2u W=6u
        MP65 N$2904 N$1046 VDD VDD p L=2u W=6u
        MN88 N$925 N$1601 GND GND n L=2u W=3u
        MN87 N$925 N$707 GND GND n L=2u W=3u
        MP93 N$924 N$916 N$921 VDD p L=2u W=3u
        MP92 N$924 N$9 N$923 VDD p L=2u W=3u
        MP91 N$923 N$1601 N$922 VDD p L=2u W=3u
        MP161 N$3696 N$3689 N$3693 VDD p L=2u W=3u
        MP160 N$3696 N$3460 N$3695 VDD p L=2u W=3u
        MP159 N$3695 N$3456 N$3694 VDD p L=2u W=3u
        MP158 N$3694 N$1017 N$3693 VDD p L=2u W=3u
        MN68 N$2908 N$1049 GND GND n L=2u W=6u
        MP23 N$28 N$2017 VDD VDD p L=2u W=3u
        MP22 N$28 N$2905 VDD VDD p L=2u W=3u
        MN27 N$31 C1 N$33 GND n L=2u W=3u
        MN26 N$31 N$24 N$32 GND n L=2u W=3u
        MN25 N$34 N$2017 GND GND n L=2u W=3u
        MN24 N$33 N$2905 N$34 GND n L=2u W=3u
        MN23 N$32 C1 GND GND n L=2u W=3u
        MN22 N$32 N$2017 GND GND n L=2u W=3u
        MP107 N$938 N$932 N$935 VDD p L=2u W=3u
        MP106 N$938 N$25 N$937 VDD p L=2u W=3u
        MP105 N$937 N$51 N$936 VDD p L=2u W=3u
        MP198 N$1020 N$1607 VDD VDD p L=2u W=3u
        MP197 N$1020 N$946 VDD VDD p L=2u W=3u
        MP196 N$1017 N$1016 VDD VDD p L=2u W=3u
        MN94 N$928 N$924 GND GND n L=2u W=3u
        MP94 N$928 N$924 VDD VDD p L=2u W=3u
        MN14 N$2020 N$15 GND GND n L=2u W=3u
        MP14 N$2020 N$15 VDD VDD p L=2u W=3u
        MP119 N$951 N$2908 N$950 VDD p L=2u W=3u
        MN260 N$4340 CLK GND GND n L=2u W=5u
        MP260 N$4340 CLK VDD VDD p L=2u W=5u
        MN259 N$4338 N$4335 GND GND n L=2u W=6u
        MP259 N$4338 N$4335 VDD VDD p L=2u W=6u
        MN258 P2 N$4338 GND GND n L=2u W=6u
        MP258 P2 N$4338 VDD VDD p L=2u W=6u
        MP257 N$4335 CLK P2 VDD p L=2u W=6u
        MN257 P2 N$4340 N$4335 GND n L=2u W=6u
        MP256 N$4336 N$4340 N$4335 VDD p L=2u W=6u
        MN256 N$4335 CLK N$4336 GND n L=2u W=6u
        MN255 N$4336 N$4339 GND GND n L=2u W=6u
        MP255 N$4336 N$4339 VDD VDD p L=2u W=6u
        MN254 N$4339 N$4337 GND GND n L=2u W=6u
        MP221 N$4324 N$4328 N$4323 VDD p L=2u W=6u
        MN221 N$4323 CLK N$4324 GND n L=2u W=6u
        MN220 N$4324 N$4327 GND GND n L=2u W=6u
        MP220 N$4324 N$4327 VDD VDD p L=2u W=6u
        MN219 N$4327 N$4325 GND GND n L=2u W=6u
        MP219 N$4327 N$4325 VDD VDD p L=2u W=6u
        MP218 N$4325 N$4328 N$4324 VDD p L=2u W=6u
        MN218 N$4324 CLK N$4325 GND n L=2u W=6u
        MP217 N$37 CLK N$4325 VDD p L=2u W=6u
        MN217 N$4325 N$4328 N$37 GND n L=2u W=6u
        MP143 N$1057 B2 VDD VDD p L=2u W=6u
        MN142 N$707 N$1055 GND GND n L=2u W=6u
        MP142 N$707 N$1055 VDD VDD p L=2u W=6u
        MP76 N$1034 A0 VDD VDD p L=2u W=6u
        MN75 N$1034 A0 N$1030 GND n L=2u W=6u
        MP75 N$1034 B2 VDD VDD p L=2u W=6u
        MN74 N$37 N$1032 GND GND n L=2u W=6u
        MP74 N$37 N$1032 VDD VDD p L=2u W=6u
        MN276 P4 N$4352 GND GND n L=2u W=6u
        MP276 P4 N$4352 VDD VDD p L=2u W=6u
        MP275 N$4349 CLK P4 VDD p L=2u W=6u
        MN275 P4 N$4354 N$4349 GND n L=2u W=6u
        MP274 N$4350 N$4354 N$4349 VDD p L=2u W=6u
        MN274 N$4349 CLK N$4350 GND n L=2u W=6u
        MN273 N$4350 N$4353 GND GND n L=2u W=6u
        MP273 N$4350 N$4353 VDD VDD p L=2u W=6u
        MN272 N$4353 N$4351 GND GND n L=2u W=6u
        MP272 N$4353 N$4351 VDD VDD p L=2u W=6u
        MP271 N$4351 N$4354 N$4350 VDD p L=2u W=6u
        MN271 N$4350 CLK N$4351 GND n L=2u W=6u
        MP270 N$4320 CLK N$4351 VDD p L=2u W=6u
        MN113 N$947 N$2908 GND GND n L=2u W=3u
        MN112 N$948 N$2908 GND GND n L=2u W=3u
        MN111 N$945 N$41 N$947 GND n L=2u W=3u
        MN110 N$947 N$1579 GND GND n L=2u W=3u
        MN109 N$946 N$945 GND GND n L=2u W=3u
        MP113 N$945 N$1579 N$944 VDD p L=2u W=3u
        MP112 N$945 N$41 N$943 VDD p L=2u W=3u
        MP111 N$944 N$2908 N$943 VDD p L=2u W=3u
        MP110 N$943 N$2908 VDD VDD p L=2u W=3u
        MP109 N$943 N$1579 VDD VDD p L=2u W=3u
        MN114 N$945 N$1579 N$948 GND n L=2u W=3u
        MP114 N$946 N$945 VDD VDD p L=2u W=3u
        MP115 N$949 N$41 VDD VDD p L=2u W=3u
        MN263 N$4346 N$4344 GND GND n L=2u W=6u
        MP263 N$4346 N$4344 VDD VDD p L=2u W=6u
        MP262 N$4344 N$4347 N$4343 VDD p L=2u W=6u
        MN262 N$4343 CLK N$4344 GND n L=2u W=6u
        MP261 N$999 CLK N$4344 VDD p L=2u W=6u
        MN261 N$4344 N$4347 N$999 GND n L=2u W=6u
        MP292 N$4362 N$4366 N$4361 VDD p L=2u W=6u
        MN292 N$4361 CLK N$4362 GND n L=2u W=6u
        MN291 N$4362 N$4365 GND GND n L=2u W=6u
        MP291 N$4362 N$4365 VDD VDD p L=2u W=6u
        MN290 N$4365 N$4363 GND GND n L=2u W=6u
        MP290 N$4365 N$4363 VDD VDD p L=2u W=6u
        MP289 N$4363 N$4366 N$4362 VDD p L=2u W=6u
        MN289 N$4362 CLK N$4363 GND n L=2u W=6u
        MP288 N$4321 CLK N$4363 VDD p L=2u W=6u
        MN288 N$4363 N$4366 N$4321 GND n L=2u W=6u
        MN287 N$4360 CLK GND GND n L=2u W=5u
        MP287 N$4360 CLK VDD VDD p L=2u W=5u
        MN286 N$4358 N$4355 GND GND n L=2u W=6u
        MP254 N$4339 N$4337 VDD VDD p L=2u W=6u
        MP253 N$4337 N$4340 N$4336 VDD p L=2u W=6u
        MN253 N$4336 CLK N$4337 GND n L=2u W=6u
        MP252 N$928 CLK N$4337 VDD p L=2u W=6u
        MN252 N$4337 N$4340 N$928 GND n L=2u W=6u
        MN251 N$4334 CLK GND GND n L=2u W=5u
        MP251 N$4334 CLK VDD VDD p L=2u W=5u
        MN250 N$4332 N$4329 GND GND n L=2u W=6u
        MP250 N$4332 N$4329 VDD VDD p L=2u W=6u
        MN249 P1 N$4332 GND GND n L=2u W=6u
        MP249 P1 N$4332 VDD VDD p L=2u W=6u
        MP248 N$4329 CLK P1 VDD p L=2u W=6u
        MN248 P1 N$4334 N$4329 GND n L=2u W=6u
        MP279 N$3704 CLK N$4357 VDD p L=2u W=6u
        MN279 N$4357 N$4360 N$3704 GND n L=2u W=6u
        MN278 N$4354 CLK GND GND n L=2u W=5u
        MP278 N$4354 CLK VDD VDD p L=2u W=5u
        MN277 N$4352 N$4349 GND GND n L=2u W=6u
        MP277 N$4352 N$4349 VDD VDD p L=2u W=6u
        MN270 N$4351 N$4354 N$4320 GND n L=2u W=6u
        MN269 N$4347 CLK GND GND n L=2u W=5u
        MP269 N$4347 CLK VDD VDD p L=2u W=5u
        MN268 N$4345 N$4342 GND GND n L=2u W=6u
        MP268 N$4345 N$4342 VDD VDD p L=2u W=6u
        MN267 P3 N$4345 GND GND n L=2u W=6u
        MP267 P3 N$4345 VDD VDD p L=2u W=6u
        MP266 N$4342 CLK P3 VDD p L=2u W=6u
        MN266 P3 N$4347 N$4342 GND n L=2u W=6u
        MP265 N$4343 N$4347 N$4342 VDD p L=2u W=6u
        MN265 N$4342 CLK N$4343 GND n L=2u W=6u
        MN264 N$4343 N$4346 GND GND n L=2u W=6u
        MP264 N$4343 N$4346 VDD VDD p L=2u W=6u
        MN295 N$4364 N$4361 GND GND n L=2u W=6u
        MP295 N$4364 N$4361 VDD VDD p L=2u W=6u
        MN294 P6 N$4364 GND GND n L=2u W=6u
        MP294 P6 N$4364 VDD VDD p L=2u W=6u
        MP293 N$4361 CLK P6 VDD p L=2u W=6u
        MN293 P6 N$4366 N$4361 GND n L=2u W=6u
        MN36 N$48 N$2906 GND GND n L=2u W=3u
        MN35 N$48 N$2904 GND GND n L=2u W=3u
        MP41 N$47 N$40 N$44 VDD p L=2u W=3u
        MN37 N$48 C1 GND GND n L=2u W=3u
        MN38 N$49 N$2904 N$50 GND n L=2u W=3u
        MP34 N$41 N$40 VDD VDD p L=2u W=3u
        MP35 N$44 C1 VDD VDD p L=2u W=3u
        MP36 N$44 N$2904 VDD VDD p L=2u W=3u
        MP136 N$3704 N$3683 VDD VDD p L=2u W=3u
        MN136 N$3704 N$3683 GND GND n L=2u W=3u
        MP149 N$3687 N$1017 VDD VDD p L=2u W=3u
        MP150 N$3687 N$3456 VDD VDD p L=2u W=3u
        MP151 N$3688 N$3456 N$3687 VDD p L=2u W=3u
        MP152 N$3689 N$3460 N$3687 VDD p L=2u W=3u
        MP195 N$1016 N$1607 N$1015 VDD p L=2u W=3u
        MP193 N$1015 N$1584 N$1014 VDD p L=2u W=3u
        MP194 N$1016 N$946 N$1014 VDD p L=2u W=3u
        MP191 N$1014 N$1607 VDD VDD p L=2u W=3u
        MP192 N$1014 N$1584 VDD VDD p L=2u W=3u
        MP6 N$9 N$6 VDD VDD p L=2u W=3u
        MN6 N$6 N$4109 N$11 GND n L=2u W=3u
        MN5 N$10 N$2907 GND GND n L=2u W=3u
        MN4 N$11 N$2907 GND GND n L=2u W=3u
        MP79 N$1035 A0 VDD VDD p L=2u W=6u
        MN78 N$1035 A0 N$1031 GND n L=2u W=6u
        MP78 N$1035 B3 VDD VDD p L=2u W=6u
        MN77 N$2017 N$1034 GND GND n L=2u W=6u
        MN62 N$4109 N$1043 GND GND n L=2u W=6u
        MP62 N$4109 N$1043 VDD VDD p L=2u W=6u
        MP68 N$2908 N$1049 VDD VDD p L=2u W=6u
        MN305 N$4372 CLK GND GND n L=2u W=5u
        MP305 N$4372 CLK VDD VDD p L=2u W=5u
        MN304 N$4370 N$4367 GND GND n L=2u W=6u
        MP304 N$4370 N$4367 VDD VDD p L=2u W=6u
        MN303 P7 N$4370 GND GND n L=2u W=6u
        MP303 P7 N$4370 VDD VDD p L=2u W=6u
        MP302 N$4367 CLK P7 VDD p L=2u W=6u
        MN302 P7 N$4372 N$4367 GND n L=2u W=6u
        MP301 N$4368 N$4372 N$4367 VDD p L=2u W=6u
        MN67 N$1050 B3 GND GND n L=2u W=6u
        MP67 N$1049 A1 VDD VDD p L=2u W=6u
        MN66 N$1049 A1 N$1050 GND n L=2u W=6u
        MN280 N$4356 CLK N$4357 GND n L=2u W=6u
        MP155 N$3693 N$3460 VDD VDD p L=2u W=3u
        MP154 N$3690 N$3689 VDD VDD p L=2u W=3u
        MN154 N$3689 N$1017 N$3692 GND n L=2u W=3u
        MN153 N$3691 N$3456 GND GND n L=2u W=3u
        MN152 N$3692 N$3456 GND GND n L=2u W=3u
        MN151 N$3689 N$3460 N$3691 GND n L=2u W=3u
        MN150 N$3691 N$1017 GND GND n L=2u W=3u
        MN149 N$3690 N$3689 GND GND n L=2u W=3u
        MP153 N$3689 N$1017 N$3688 VDD p L=2u W=3u
        MP156 N$3693 N$1017 VDD VDD p L=2u W=3u
        MN186 N$1011 N$2902 N$1012 GND n L=2u W=3u
        MN185 N$1010 N$2494 GND GND n L=2u W=3u
        MN184 N$1010 N$956 GND GND n L=2u W=3u
        MN190 N$3451 N$1009 GND GND n L=2u W=3u
        MP190 N$3451 N$1009 VDD VDD p L=2u W=3u
        MN165 N$988 N$2903 N$990 GND n L=2u W=3u
        MN189 N$1009 N$2494 N$1011 GND n L=2u W=3u
        MN192 N$1018 N$1607 GND GND n L=2u W=3u
        MN193 N$1016 N$946 N$1018 GND n L=2u W=3u
        MN188 N$1009 N$1002 N$1010 GND n L=2u W=3u
        MN162 N$4321 N$3696 GND GND n L=2u W=3u
        MP162 N$4321 N$3696 VDD VDD p L=2u W=3u
        MN161 N$3696 N$3460 N$3698 GND n L=2u W=3u
        MN160 N$3696 N$3689 N$3697 GND n L=2u W=3u
        MN159 N$3699 N$3456 GND GND n L=2u W=3u
        MN158 N$3698 N$1017 N$3699 GND n L=2u W=3u
        MN157 N$3697 N$3460 GND GND n L=2u W=3u
        MN156 N$3697 N$3456 GND GND n L=2u W=3u
        MN155 N$3697 N$1017 GND GND n L=2u W=3u
        MN187 N$1012 N$956 GND GND n L=2u W=3u
        MN205 N$1077 A3 N$1062 GND n L=2u W=6u
        MP205 N$1077 B1 VDD VDD p L=2u W=6u
        MN104 N$940 N$1578 N$941 GND n L=2u W=3u
        MN148 N$1584 N$1059 GND GND n L=2u W=6u
        MP148 N$1584 N$1059 VDD VDD p L=2u W=6u
        MN147 N$1060 B3 GND GND n L=2u W=6u
        MP147 N$1059 A2 VDD VDD p L=2u W=6u
        MN146 N$1059 A2 N$1060 GND n L=2u W=6u
        MP146 N$1059 B3 VDD VDD p L=2u W=6u
        MN145 N$1579 N$1057 GND GND n L=2u W=6u
        MP145 N$1579 N$1057 VDD VDD p L=2u W=6u
        MP206 N$1077 A3 VDD VDD p L=2u W=6u
        MN137 N$1051 A2 N$1053 GND n L=2u W=6u
        MP137 N$1051 B1 VDD VDD p L=2u W=6u
        MP139 N$1578 N$1051 VDD VDD p L=2u W=6u
        MN138 N$1053 B1 GND GND n L=2u W=6u
        MP71 N$2907 N$1033 VDD VDD p L=2u W=6u
        MN70 N$1029 B1 GND GND n L=2u W=6u
        MP70 N$1033 A0 VDD VDD p L=2u W=6u
        MN69 N$1033 A0 N$1029 GND n L=2u W=6u
        MP69 N$1033 B1 VDD VDD p L=2u W=6u
        MN143 N$1057 A2 N$1058 GND n L=2u W=6u
        MP213 N$1607 N$1066 VDD VDD p L=2u W=6u
        MN216 N$3456 N$1068 GND GND n L=2u W=6u
        MP216 N$3456 N$1068 VDD VDD p L=2u W=6u
        MP247 N$4330 N$4334 N$4329 VDD p L=2u W=6u
        MN247 N$4329 CLK N$4330 GND n L=2u W=6u
        MN246 N$4330 N$4333 GND GND n L=2u W=6u
        MP246 N$4330 N$4333 VDD VDD p L=2u W=6u
        MN245 N$4333 N$4331 GND GND n L=2u W=6u
        MP245 N$4333 N$4331 VDD VDD p L=2u W=6u
        MN49 N$3671 N$3451 GND GND n L=2u W=3u
        MN50 N$3671 N$3701 GND GND n L=2u W=3u
        MN51 N$3671 C1 GND GND n L=2u W=3u
        MN52 N$3672 N$3451 N$3673 GND n L=2u W=3u
        MN48 N$3664 N$3451 N$3666 GND n L=2u W=3u
        MP48 N$3700 N$3664 VDD VDD p L=2u W=3u
        MP49 N$3667 C1 VDD VDD p L=2u W=3u
        MP50 N$3667 N$3451 VDD VDD p L=2u W=3u
        MP51 N$3667 N$3701 VDD VDD p L=2u W=3u
        MP52 N$3668 N$3451 N$3667 VDD p L=2u W=3u
        MP53 N$3669 N$3701 N$3668 VDD p L=2u W=3u
        MP55 N$3670 N$3664 N$3667 VDD p L=2u W=3u
        MP54 N$3670 C1 N$3669 VDD p L=2u W=3u
        MN176 N$999 N$995 GND GND n L=2u W=3u
        MN47 N$3665 N$3701 GND GND n L=2u W=3u
        MN80 N$2906 N$1035 GND GND n L=2u W=6u
        MP80 N$2906 N$1035 VDD VDD p L=2u W=6u
        MN79 N$1031 B3 GND GND n L=2u W=6u
        MN61 N$1044 B0 GND GND n L=2u W=6u
        MP61 N$1043 A1 VDD VDD p L=2u W=6u
        MN60 N$1043 A1 N$1044 GND n L=2u W=6u
        MP60 N$1043 B0 VDD VDD p L=2u W=6u
        MN59 N$2905 N$1038 GND GND n L=2u W=6u
        MP59 N$2905 N$1038 VDD VDD p L=2u W=6u
        MN58 N$1041 B1 GND GND n L=2u W=6u
        MN64 N$1047 B2 GND GND n L=2u W=6u
        MP64 N$1046 A1 VDD VDD p L=2u W=6u
        MN63 N$1046 A1 N$1047 GND n L=2u W=6u
        MP63 N$1046 B2 VDD VDD p L=2u W=6u
        MP3 N$5 N$2907 N$2 VDD p L=2u W=3u
        MP2 N$2 N$2907 VDD VDD p L=2u W=3u
        MP1 N$2 N$4109 VDD VDD p L=2u W=3u
        MP77 N$2017 N$1034 VDD VDD p L=2u W=6u
        MN57 N$1038 A1 N$1041 GND n L=2u W=6u
        MN141 N$1056 B0 GND GND n L=2u W=6u
        MP57 N$1038 B1 VDD VDD p L=2u W=6u
        MP58 N$1038 A1 VDD VDD p L=2u W=6u
        MN76 N$1030 B2 GND GND n L=2u W=6u
        MN55 N$3670 C1 N$3672 GND n L=2u W=3u
        MN54 N$3670 N$3664 N$3671 GND n L=2u W=3u
        MN53 N$3673 N$3701 GND GND n L=2u W=3u

*.ends mynand3

* Auxiliary circuit for power analysis
Cp Pav 0 100p
Rp Pav 0 100k
Fp 0 Pav Vtstp 0.003125
*Output load capacitance if you have any

*Cload1 out GND 200fF
.MODEL n NMOS LEVEL = 3
+ TOX = 200E-10 NSUB = 1E17 GAMMA = 0.5
+ PHI = 0.7 VTO = 0.8 DELTA = 3.0
+ UO = 650 ETA = 3.0E-6 THETA = 0.1
+ KP = 120E-6 VMAX = 1E5 KAPPA = 0.3
+ RSH = 0 NFS = 1E12 TPG = 1
+ XJ = 500E-9 LD = 100E-9
+ CGDO = 200E-12 CGSO = 200E-12 CGBO = 1E-10
+ CJ = 400E-6 PB = 1 MJ = 0.5
+ CJSW = 300E-12 MJSW = 0.5

.MODEL p PMOS LEVEL = 3
+ TOX = 200E-10 NSUB = 1E17 GAMMA = 0.6
+ PHI = 0.7 VTO = -0.9 DELTA = 0.1
+ UO = 250 ETA = 0 THETA = 0.1
+ KP = 40E-6 VMAX = 5E4 KAPPA = 1
+ RSH = 0 NFS = 1E12 TPG = -1
+ XJ = 500E-9 LD = 100E-9
+ CGDO = 200E-12 CGSO = 200E-12 CGBO = 1E-10
+ CJ = 400E-6 PB = 1 MJ = 0.5
+ CJSW = 300E-12 MJSW = 0.5

*Define power rails
Vddt top 0 5
Vtstp top Vdd 0
Vss GND 0 0

* Define input voltages of A and B

Vclk CLK 0 PWL(0 5 20N 5 20.1N 0 40N 0 40.1N 5 60N 5 60.1N 0 80N 0 80.1N 5
+ 100N 5 100.1N 0 120N 0 120.1N 5 140N 5 140.1N 0 160N 0 160.1N 5 180N 5 180.1N 0 200N 0)
Va0 A0 0 PWL(0 5 20N 5 20.1N 5 40N 5 40.1N 5 60N 5 60.1N 5 80N 5 80.1N 5
+ 100N 5 100.1N 5 120N 5 120.1N 5 140N 5 140.1N 5 160N 5 160.1N 5 180N 5 180.1N 5 200N 5)
Va2 A2 0 PWL(0 0 20N 0 20.1N 0 40N 0 40.1N 0 60N 0 60.1N 0 80N 0 80.1N 0
+ 100N 0 100.1N 0 120N 0 120.1N 0 140N 0 140.1N 0 160N 0 160.1N 0 180N 0 180.1N 0 200N 0)
Va1 A1 0 PWL(0 5 20N 5 20.1N 5 40N 5 40.1N 5 60N 5 60.1N 5 80N 5 80.1N 5
+ 100N 5 100.1N 5 120N 5 120.1N 5 140N 5 140.1N 5 160N 5 160.1N 5 180N 5 180.1N 5 200N 5)
Va3 A3 0 PWL(0 0 20N 0 20.1N 0 40N 0 40.1N 0 60N 0 60.1N 0 80N 0 80.1N 0
+ 100N 0 100.1N 0 120N 0 120.1N 0 140N 0 140.1N 0 160N 0 160.1N 0 180N 0 180.1N 0 200N 0)
Vrst1 RST1 0 PWL(0 5 20N 5 20.1N 5 40N 5 40.1N 0 60N 0 60.1N 0 80N 0 80.1N 0
+ 100N 0 100.1N 0 120N 0 120.1N 0 140N 0 140.1N 0 160N 0 160.1N 0 180N 0 180.1N 0 200N 0)
Vb0 B0 0 PWL(0 5 20N 5 20.1N 5 40N 5 40.1N 5 60N 5 60.1N 5 80N 5 80.1N 5
+ 100N 5 100.1N 5 120N 5 120.1N 5 140N 5 140.1N 5 160N 5 160.1N 5 180N 5 180.1N 5 200N 5)
Vb2 B2 0 PWL(0 0 20N 0 20.1N 0 40N 0 40.1N 0 60N 0 60.1N 0 80N 0 80.1N 0
+ 100N 0 100.1N 0 120N 0 120.1N 0 140N 0 140.1N 0 160N 0 160.1N 0 180N 0 180.1N 0 200N 0)
Vb1 B1 0 PWL(0 5 20N 5 20.1N 5 40N 5 40.1N 5 60N 5 60.1N 5 80N 5 80.1N 5
+ 100N 5 100.1N 5 120N 5 120.1N 5 140N 5 140.1N 5 160N 5 160.1N 5 180N 5 180.1N 5 200N 5)
Vb3 B3 0 PWL(0 0 20N 0 20.1N 0 40N 0 40.1N 0 60N 0 60.1N 0 80N 0 80.1N 0
+ 100N 0 100.1N 0 120N 0 120.1N 0 140N 0 140.1N 0 160N 0 160.1N 0 180N 0 180.1N 0 200N 0)
Vc1 C1 0 PWL(0 0 20N 0 20.1N 0 40N 0 40.1N 0 60N 0 60.1N 0 80N 0 80.1N 0
+ 100N 0 100.1N 0 120N 0 120.1N 0 140N 0 140.1N 0 160N 0 160.1N 0 180N 0 180.1N 0 200N 0)



*Define transient simulation and probe voltage/current signals
.TRAN 20N 200N
.PROBE V(*) I(*)
.end