*
* .CONNECT statements
*
.CONNECT GND 0


* ELDO netlist generated with ICnet by 'mentor' on Mon Mar 17 2008 at 15:04:13

*
* Globals.
*
.global VDD GND

*
* MAIN CELL: Component pathname : /home/mentor/EXOR/exor
*
        MN6 N$11 B GND GND n L=2u W=6u
        MP6 N$11 B VDD VDD p L=2u W=6u
        MN5 N$5 A GND GND n L=2u W=6u
        MP5 N$5 A VDD VDD p L=2u W=6u
        MN4 N$8 N$11 GND GND n L=2u W=6u
        MN3 OUT A N$8 GND n L=2u W=6u
        MN2 N$6 B GND GND n L=2u W=6u
        MN1 OUT N$5 N$6 GND n L=2u W=6u
        MP4 OUT B N$4 VDD p L=2u W=6u
        MP3 N$4 N$11 VDD VDD p L=2u W=6u
        MP2 OUT N$5 N$4 VDD p L=2u W=6u
        MP1 N$4 A VDD VDD p L=2u W=6u
*
.end
