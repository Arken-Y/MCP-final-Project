




*.subckt mynand3 A B GND Out Vdd



* MAIN CELL: Component pathname : /home/mentor/jack/jaggu
*
               MN71 N$66 N$65 GND GND n L=2u W=5u
        MN77 N$72 N$71 GND GND n L=2u W=5u
        MP77 N$72 N$71 VDD VDD p L=2u W=5u
        MN76 N$71 N$61 GND GND n L=2u W=5u
        MN75 N$71 N$60 GND GND n L=2u W=5u
        MP76 N$71 N$61 N$70 VDD p L=2u W=5u
        MP75 N$70 N$60 VDD VDD p L=2u W=5u
        MN80 N$75 N$74 GND GND n L=2u W=5u
        MP80 N$75 N$74 VDD VDD p L=2u W=5u
        MN79 N$74 N$63 GND GND n L=2u W=5u
        MN78 N$74 N$62 GND GND n L=2u W=5u
        MP79 N$74 N$63 N$73 VDD p L=2u W=5u
        MP78 N$73 N$62 VDD VDD p L=2u W=5u
        MN951 N$14074 N$11345 GND GND n L=2u W=5u
        MP951 N$14074 N$11345 VDD VDD p L=2u W=5u
        MN950 N$14078 N$14074 N$66 GND n L=2u W=5u
        MP950 N$66 N$11345 N$14078 VDD p L=2u W=5u
        MN949 N$14078 N$11345 GND GND n L=2u W=5u
        MP949 GND N$14074 N$14078 VDD p L=2u W=5u
        MP957 N$75 N$11345 N$14081 VDD p L=2u W=5u
        MN956 N$14081 N$11345 GND GND n L=2u W=5u
        MP956 GND N$14074 N$14081 VDD p L=2u W=5u
        MN955 N$14080 N$14074 N$72 GND n L=2u W=5u
        MP955 N$72 N$11345 N$14080 VDD p L=2u W=5u
        MN954 N$14080 N$11345 GND GND n L=2u W=5u
        MP954 GND N$14074 N$14080 VDD p L=2u W=5u
        MN953 N$14079 N$14074 N$415 GND n L=2u W=5u
        MP953 N$415 N$11345 N$14079 VDD p L=2u W=5u
        MN952 N$14079 N$11345 GND GND n L=2u W=5u
        MP952 GND N$14074 N$14079 VDD p L=2u W=5u
        MN957 N$14081 N$14074 N$75 GND n L=2u W=5u
        MN53 N$14093 N$420 N$60 GND n L=2u W=6u
        MP53 N$14093 N$417 N$60 VDD p L=2u W=6u
        MP52 GND N$421 N$59 VDD p L=2u W=6u
        MN52 GND N$419 N$59 GND n L=2u W=6u
        MN51 N$36 N$421 N$59 GND n L=2u W=6u
        MP51 N$36 N$419 N$59 VDD p L=2u W=6u
        MP50 GND N$420 N$58 VDD p L=2u W=6u
        MP57 N$14092 N$417 N$62 VDD p L=2u W=6u
        MP56 GND N$421 N$61 VDD p L=2u W=6u
        MN56 GND N$419 N$61 GND n L=2u W=6u
        MN55 N$25 N$421 N$61 GND n L=2u W=6u
        MP55 N$25 N$419 N$61 VDD p L=2u W=6u
        MP54 GND N$420 N$60 VDD p L=2u W=6u
        MN60 GND N$419 N$63 GND n L=2u W=6u
        MN59 N$46 N$421 N$63 GND n L=2u W=6u
        MP59 N$46 N$419 N$63 VDD p L=2u W=6u
        MP58 GND N$420 N$62 VDD p L=2u W=6u
        MN58 GND N$417 N$62 GND n L=2u W=6u
        MN57 N$14092 N$420 N$62 GND n L=2u W=6u
        MP71 N$66 N$65 VDD VDD p L=2u W=5u
        MN70 N$65 N$56 GND GND n L=2u W=5u
        MN69 N$65 N$53 GND GND n L=2u W=5u
        MP70 N$65 N$56 N$64 VDD p L=2u W=5u
        MP69 N$64 N$53 VDD VDD p L=2u W=5u
        MP60 GND N$421 N$63 VDD p L=2u W=6u
        MN74 N$415 N$68 GND GND n L=2u W=5u
        MP74 N$415 N$68 VDD VDD p L=2u W=5u
        MN73 N$68 N$59 GND GND n L=2u W=5u
        MN72 N$68 N$58 GND GND n L=2u W=5u
        MP73 N$68 N$59 N$67 VDD p L=2u W=5u
        MP72 N$67 N$58 VDD VDD p L=2u W=5u
        MN37 N$42 N$38 GND GND n L=2u W=6u
        MP37 N$42 N$38 VDD VDD p L=2u W=6u
        MN36 N$45 N$43 GND GND n L=2u W=6u
        MN35 N$41 N$38 N$45 GND n L=2u W=6u
        MN34 N$44 N$26 GND GND n L=2u W=6u
        MN33 N$41 N$42 N$44 GND n L=2u W=6u
        MP41 N$28 N$14045 VDD VDD p L=2u W=6u
        MN40 H_A_COUT N$37 GND GND n L=2u W=6u
        MP40 H_A_COUT N$37 VDD VDD p L=2u W=6u
        MN39 N$46 N$41 GND GND n L=2u W=6u
        MP39 N$46 N$41 VDD VDD p L=2u W=6u
        MN38 N$43 N$26 GND GND n L=2u W=6u
        MP44 N$16 N$14093 VDD VDD p L=2u W=6u
        MN43 N$3 N$14046 GND GND n L=2u W=6u
        MP43 N$3 N$14046 VDD VDD p L=2u W=6u
        MN42 N$38 N$14092 GND GND n L=2u W=6u
        MP42 N$38 N$14092 VDD VDD p L=2u W=6u
        MN41 N$28 N$14045 GND GND n L=2u W=6u
        MN47 N$13 N$421 N$56 GND n L=2u W=6u
        MP47 N$13 N$419 N$56 VDD p L=2u W=6u
        MP46 GND N$420 N$53 VDD p L=2u W=6u
        MN46 GND N$417 N$53 GND n L=2u W=6u
        MN45 N$14046 N$420 N$53 GND n L=2u W=6u
        MP45 N$14046 N$417 N$53 VDD p L=2u W=6u
        MN44 N$16 N$14093 GND GND n L=2u W=6u
        MN50 GND N$417 N$58 GND n L=2u W=6u
        MN49 N$14045 N$420 N$58 GND n L=2u W=6u
        MP49 N$14045 N$417 N$58 VDD p L=2u W=6u
        MP48 GND N$421 N$56 VDD p L=2u W=6u
        MN48 GND N$419 N$56 GND n L=2u W=6u
        MN54 GND N$417 N$60 GND n L=2u W=6u
        MP22 N$27 N$14 VDD VDD p L=2u W=6u
        MP21 N$27 N$28 VDD VDD p L=2u W=6u
        MN20 N$26 N$15 GND GND n L=2u W=6u
        MP20 N$26 N$15 VDD VDD p L=2u W=6u
        MN19 N$25 N$20 GND GND n L=2u W=6u
        MN23 N$31 N$32 N$34 GND n L=2u W=6u
        MP26 N$31 N$14 N$30 VDD p L=2u W=6u
        MP25 N$30 N$33 VDD VDD p L=2u W=6u
        MP24 N$31 N$32 N$30 VDD p L=2u W=6u
        MP23 N$30 N$28 VDD VDD p L=2u W=6u
        MN22 N$29 N$28 GND GND n L=2u W=6u
        MN28 N$33 N$14 GND GND n L=2u W=6u
        MP28 N$33 N$14 VDD VDD p L=2u W=6u
        MN27 N$32 N$28 GND GND n L=2u W=6u
        MP27 N$32 N$28 VDD VDD p L=2u W=6u
        MN26 N$35 N$33 GND GND n L=2u W=6u
        MN25 N$31 N$28 N$35 GND n L=2u W=6u
        MN24 N$34 N$14 GND GND n L=2u W=6u
        MP32 N$37 N$26 VDD VDD p L=2u W=6u
        MP31 N$37 N$38 VDD VDD p L=2u W=6u
        MN30 N$17 N$27 GND GND n L=2u W=6u
        MP30 N$17 N$27 VDD VDD p L=2u W=6u
        MN29 N$36 N$31 GND GND n L=2u W=6u
        MP29 N$36 N$31 VDD VDD p L=2u W=6u
        MP36 N$41 N$26 N$40 VDD p L=2u W=6u
        MP35 N$40 N$43 VDD VDD p L=2u W=6u
        MP34 N$41 N$42 N$40 VDD p L=2u W=6u
        MP33 N$40 N$38 VDD VDD p L=2u W=6u
        MN32 N$39 N$38 GND GND n L=2u W=6u
        MN31 N$37 N$26 N$39 GND n L=2u W=6u
        MP38 N$43 N$26 VDD VDD p L=2u W=6u
        MP324 GND N$348 N$14087 VDD p L=2u W=5u
        MP325 N$317 N$11347 N$14087 VDD p L=2u W=5u
        MN740 N$11088 N$11327 N$11330 GND n L=2u W=6u
        MP739 N$11328 N$11327 N$11330 VDD p L=2u W=6u
        MN739 N$11330 CK N$11328 GND n L=2u W=6u
        MN738 N$11328 N$11329 GND GND n L=2u W=6u
        MN767 N$11347 N$11345 GND GND n L=2u W=5u
        MP767 N$11347 N$11345 VDD VDD p L=2u W=5u
        MN766 N$11345 N$11088 GND GND n L=2u W=5u
        MN747 N$11345 N$11344 GND GND n L=2u W=5u
        MN365 N$390 N$409 N$376 GND n L=2u W=5u
        MP365 N$376 N$14096 N$390 VDD p L=2u W=5u
        MN364 N$390 N$14096 GND GND n L=2u W=5u
        MP364 GND N$409 N$390 VDD p L=2u W=5u
        MN363 N$389 N$409 N$411 GND n L=2u W=5u
        MP363 N$411 N$14096 N$389 VDD p L=2u W=5u
        MN362 N$389 N$14096 P4 GND n L=2u W=5u
        MP362 P4 N$409 N$389 VDD p L=2u W=5u
        MP97 N$99 N$386 N$96 VDD p L=2u W=3u
        MP5 N$7 N$10 VDD VDD p L=2u W=6u
        MP4 N$8 N$9 N$7 VDD p L=2u W=6u
        MP3 N$7 N$3 VDD VDD p L=2u W=6u
        MP740 N$11330 CK N$11088 VDD p L=2u W=6u
        MP271 N$312 N$313 N$314 VDD p L=2u W=6u
        MN271 N$314 CK N$312 GND n L=2u W=6u
        MP270 N$250 CK N$312 VDD p L=2u W=6u
        MN270 N$312 N$313 N$250 GND n L=2u W=6u
        MN269 N$306 CK GND GND n L=2u W=5u
        MN737 N$11329 N$11326 GND GND n L=2u W=6u
        MP737 N$11329 N$11326 VDD VDD p L=2u W=6u
        MP736 N$11326 N$11327 N$11328 VDD p L=2u W=6u
        MP741 N$11088 N$11331 VDD VDD p L=2u W=6u
        MN310 N$344 CK N$342 GND n L=2u W=6u
        MN309 N$342 N$343 GND GND n L=2u W=6u
        MN350 N$397 N$11347 N$338 GND n L=2u W=5u
        MP350 N$338 N$14095 N$397 VDD p L=2u W=5u
        MN349 N$397 N$14095 N$14090 GND n L=2u W=5u
        MP338 N$296 N$14095 N$372 VDD p L=2u W=5u
        MN337 N$372 N$14095 N$14084 GND n L=2u W=5u
        MP337 N$14084 N$11347 N$372 VDD p L=2u W=5u
        MN336 N$14095 N$11347 GND GND n L=2u W=5u
        MP336 N$14095 N$11347 VDD VDD p L=2u W=5u
        MN335 N$398 N$11347 N$361 GND n L=2u W=5u
        MP335 N$361 N$14095 N$398 VDD p L=2u W=5u
        MP371 N$396 N$14096 N$395 VDD p L=2u W=5u
        MN370 N$395 N$14096 GND GND n L=2u W=5u
        MN7 N$9 N$3 GND GND n L=2u W=6u
        MP7 N$9 N$3 VDD VDD p L=2u W=6u
        MN357 N$386 N$409 N$372 GND n L=2u W=5u
        MN161 N$182 N$390 GND GND n L=2u W=3u
        MN160 N$181 N$14078 N$182 GND n L=2u W=3u
        MN159 N$180 N$156 GND GND n L=2u W=3u
        MN158 N$180 N$390 GND GND n L=2u W=3u
        MN157 N$180 N$14078 GND GND n L=2u W=3u
        MN322 N$14086 N$11347 GND GND n L=2u W=5u
        MP322 GND N$348 N$14086 VDD p L=2u W=5u
        MN321 N$14085 N$348 N$384 GND n L=2u W=5u
        MP321 N$384 N$11347 N$14085 VDD p L=2u W=5u
        MN320 N$14085 N$11347 GND GND n L=2u W=5u
        MP158 N$176 N$14078 VDD VDD p L=2u W=3u
        MP157 N$176 N$156 VDD VDD p L=2u W=3u
        MP186 N$210 N$14080 VDD VDD p L=2u W=3u
        MN717 N$11314 N$11315 N$382 GND n L=2u W=6u
        MP361 N$374 N$14096 N$388 VDD p L=2u W=5u
        MN186 N$214 N$394 GND GND n L=2u W=3u
        MN185 N$214 N$14080 GND GND n L=2u W=3u
        MP191 N$213 N$205 N$210 VDD p L=2u W=3u
        MP190 N$213 N$190 N$212 VDD p L=2u W=3u
        MP189 N$212 N$394 N$211 VDD p L=2u W=3u
        MP188 N$211 N$14080 N$210 VDD p L=2u W=3u
        MP213 N$148 N$265 N$246 VDD p L=2u W=5u
        MN10 N$14 N$2 GND GND n L=2u W=6u
        MP729 N$11322 N$11323 VDD VDD p L=2u W=6u
        MN728 N$11323 N$11320 GND GND n L=2u W=6u
        MP728 N$11323 N$11320 VDD VDD p L=2u W=6u
        MP727 N$11320 N$11321 N$11322 VDD p L=2u W=6u
        MN727 N$11322 CK N$11320 GND n L=2u W=6u
        MP726 N$14096 CK N$11320 VDD p L=2u W=6u
        MN726 N$11320 N$11321 N$14096 GND n L=2u W=6u
        MN725 N$11315 CK GND GND n L=2u W=5u
        MP725 N$11315 CK VDD VDD p L=2u W=5u
        MP82 N$77 N$385 VDD VDD p L=2u W=3u
        MP81 N$77 GND VDD VDD p L=2u W=3u
        MN83 N$81 GND N$85 GND n L=2u W=3u
        MN82 N$85 GND GND GND n L=2u W=3u
        MN81 N$84 N$81 GND GND n L=2u W=3u
        MP723 N$14096 N$11319 VDD VDD p L=2u W=6u
        MP722 N$11318 CK N$14096 VDD p L=2u W=6u
        MN722 N$14096 N$11315 N$11318 GND n L=2u W=6u
        MP747 N$11108 N$11344 N$11104 VDD p L=2u W=5u
        MP746 N$11104 N$11099 N$11100 VDD p L=2u W=5u
        MP745 N$11100 N$14096 N$11096 VDD p L=2u W=5u
        MP744 N$11096 N$382 VDD VDD p L=2u W=5u
        MP749 N$11332 N$11333 N$11334 VDD p L=2u W=6u
        MN749 N$11334 CK N$11332 GND n L=2u W=6u
        MP748 N$11083 CK N$11332 VDD p L=2u W=6u
        MN378 N$1539 N$11787 GND GND n L=2u W=6u
        MP378 N$1539 N$11787 VDD VDD p L=2u W=6u
        MP663 N$1488 N$1416 N$1521 VDD p L=2u W=5u
        MN662 N$1450 N$1485 GND GND n L=2u W=3u
        MP662 N$1450 N$1485 VDD VDD p L=2u W=3u
        MN661 N$1435 N$1484 GND GND n L=2u W=3u
        MN693 N$1398 N$1397 GND GND n L=2u W=6u
        MN694 N$1396 CK N$1398 GND n L=2u W=6u
        MN688 N$1401 N$1402 GND GND n L=2u W=6u
        MP693 N$1398 N$1397 VDD VDD p L=2u W=6u
        MP11 N$15 N$16 VDD VDD p L=2u W=6u
        MN338 N$372 N$11347 N$296 GND n L=2u W=5u
        MP383 N$11778 N$11781 VDD VDD p L=2u W=6u
        MP382 N$11781 N$11780 N$11779 VDD p L=2u W=6u
        MN382 N$11779 CK N$11781 GND n L=2u W=6u
        MP388 N$11775 N$11777 VDD VDD p L=2u W=6u
        MN387 N$12632 N$11775 GND GND n L=2u W=6u
        MP387 N$12632 N$11775 VDD VDD p L=2u W=6u
        MP386 N$11777 CK N$12632 VDD p L=2u W=6u
        MN386 N$12632 N$11780 N$11777 GND n L=2u W=6u
        MP385 N$11779 N$11780 N$11777 VDD p L=2u W=6u
        MN385 N$11777 CK N$11779 GND n L=2u W=6u
        MN372 N$11784 N$11789 N$11570 GND n L=2u W=6u
        MN176 N$196 N$188 N$197 GND n L=2u W=3u
        MN175 N$199 N$392 GND GND n L=2u W=3u
        MN342 N$374 N$11347 N$310 GND n L=2u W=5u
        MP342 N$310 N$14095 N$374 VDD p L=2u W=5u
        MN341 N$374 N$14095 N$14086 GND n L=2u W=5u
        MP341 N$14086 N$11347 N$374 VDD p L=2u W=5u
        MN188 N$215 N$14080 N$216 GND n L=2u W=3u
        MN187 N$214 N$190 GND GND n L=2u W=3u
        MN110 N$121 GND GND GND n L=2u W=3u
        MN109 N$120 N$118 GND GND n L=2u W=3u
        MN138 N$157 GND GND GND n L=2u W=3u
        MN137 N$156 N$154 GND GND n L=2u W=3u
        MP141 N$154 GND N$153 VDD p L=2u W=3u
        MP140 N$154 N$138 N$150 VDD p L=2u W=3u
        MP139 N$153 N$389 N$150 VDD p L=2u W=3u
        MN319 N$14084 N$348 N$296 GND n L=2u W=5u
        MN328 N$14088 N$348 N$324 GND n L=2u W=5u
        MP328 N$324 N$11347 N$14088 VDD p L=2u W=5u
        MN327 N$14088 N$11347 GND GND n L=2u W=5u
        MP327 GND N$348 N$14088 VDD p L=2u W=5u
        MP326 GND N$348 N$14091 VDD p L=2u W=5u
        MN332 N$14090 N$348 N$338 GND n L=2u W=5u
        MP332 N$338 N$11347 N$14090 VDD p L=2u W=5u
        MN179 N$207 N$205 GND GND n L=2u W=3u
        MP183 N$205 N$14080 N$204 VDD p L=2u W=3u
        MP182 N$205 N$190 N$202 VDD p L=2u W=3u
        MP330 N$331 N$11347 N$14089 VDD p L=2u W=5u
        MP297 N$262 CK N$333 VDD p L=2u W=6u
        MN297 N$333 N$334 N$262 GND n L=2u W=6u
        MP708 N$1408 CK N$1388 VDD p L=2u W=6u
        MN333 N$14091 N$348 N$345 GND n L=2u W=5u
        MN12 N$18 N$16 GND GND n L=2u W=6u
        MN11 N$15 N$17 N$18 GND n L=2u W=6u
        MN729 N$11322 N$11323 GND GND n L=2u W=6u
        MN730 N$11324 CK N$11322 GND n L=2u W=6u
        MP730 N$11322 N$11321 N$11324 VDD p L=2u W=6u
        MP85 N$81 GND N$80 VDD p L=2u W=3u
        MP84 N$81 GND N$77 VDD p L=2u W=3u
        MP673 GND N$1557 N$14097 VDD p L=2u W=5u
        MN672 N$14097 N$1557 N$1467 GND n L=2u W=5u
        MP15 N$19 N$22 VDD VDD p L=2u W=6u
        MP14 N$20 N$21 N$19 VDD p L=2u W=6u
        MP13 N$19 N$16 VDD VDD p L=2u W=6u
        MN97 N$100 N$84 N$103 GND n L=2u W=3u
        MN96 N$103 GND GND GND n L=2u W=3u
        MN890 N$14028 N$14040 GND GND n L=2u W=5u
        MP891 P1 N$14040 N$14027 VDD p L=2u W=5u
        MN334 N$398 N$14095 OUT8 GND n L=2u W=5u
        MP343 N$14087 N$11347 N$411 VDD p L=2u W=5u
        MN702 N$1392 N$1391 GND GND n L=2u W=6u
        MP702 N$1392 N$1391 VDD VDD p L=2u W=6u
        MN701 N$1391 N$1394 GND GND n L=2u W=6u
        MP701 N$1391 N$1394 VDD VDD p L=2u W=6u
        MP707 N$1393 CK VDD VDD p L=2u W=5u
        MN706 N$1389 N$1390 GND GND n L=2u W=6u
        MP706 N$1389 N$1390 VDD VDD p L=2u W=6u
        MN705 N$14093 N$1389 GND GND n L=2u W=6u
        MP705 N$14093 N$1389 VDD VDD p L=2u W=6u
        MP704 N$1390 CK N$14093 VDD p L=2u W=6u
        MN704 N$14093 N$1393 N$1390 GND n L=2u W=6u
        MP710 N$1385 N$1388 VDD VDD p L=2u W=6u
        MP709 N$1388 N$1387 N$1386 VDD p L=2u W=6u
        MN709 N$1386 CK N$1388 GND n L=2u W=6u
        MN296 N$327 CK GND GND n L=2u W=5u
        MP296 N$327 CK VDD VDD p L=2u W=5u
        MN84 N$86 N$385 GND GND n L=2u W=3u
        MN112 N$122 N$387 GND GND n L=2u W=3u
        MN111 N$118 N$102 N$121 GND n L=2u W=3u
        MP542 N$11813 RST VDD VDD p L=2u W=5u
        MP574 N$1507 N$1509 VDD VDD p L=2u W=6u
        MP551 N$1530 N$1539 VDD VDD p L=2u W=5u
        MN550 N$1529 N$1530 GND GND n L=2u W=5u
        MP550 GND N$1539 N$1529 VDD p L=2u W=5u
        MN549 N$1529 N$1539 N$1539 GND n L=2u W=5u
        MP549 N$1539 N$1530 N$1529 VDD p L=2u W=5u
        MP666 N$1486 N$1416 N$1512 VDD p L=2u W=5u
        MP691 N$1400 N$1399 N$1398 VDD p L=2u W=6u
        MP697 N$1395 N$1396 VDD VDD p L=2u W=6u
        MN696 N$14045 N$1395 GND GND n L=2u W=6u
        MP696 N$14045 N$1395 VDD VDD p L=2u W=6u
        MP695 N$1396 CK N$14045 VDD p L=2u W=6u
        MN695 N$14045 N$1399 N$1396 GND n L=2u W=6u
        MP694 N$1398 N$1399 N$1396 VDD p L=2u W=6u
        MP700 N$1394 N$1393 N$1392 VDD p L=2u W=6u
        MP659 N$1481 N$1488 VDD VDD p L=2u W=3u
        MN659 N$1481 N$1488 GND GND n L=2u W=3u
        MP660 N$1465 N$1486 VDD VDD p L=2u W=3u
        MN658 N$1422 N$1426 GND GND n L=2u W=3u
        MN697 N$1395 N$1396 GND GND n L=2u W=6u
        MP703 N$1392 N$1393 N$1390 VDD p L=2u W=6u
        MN703 N$1390 CK N$1392 GND n L=2u W=6u
        MP670 N$1484 N$1416 N$1496 VDD p L=2u W=5u
        MN669 N$1504 N$1416 N$1526 GND n L=2u W=5u
        MP675 N$1452 N$1413 N$1410 VDD p L=2u W=5u
        MN674 N$1413 N$1557 GND GND n L=2u W=5u
        MP674 N$1413 N$1557 VDD VDD p L=2u W=5u
        MN673 N$14097 N$1413 GND GND n L=2u W=5u
        MN759 N$11341 N$11338 GND GND n L=2u W=6u
        MP759 N$11341 N$11338 VDD VDD p L=2u W=6u
        MP758 N$11338 N$11339 N$11340 VDD p L=2u W=6u
        MN758 N$11340 CK N$11338 GND n L=2u W=6u
        MP757 N$11099 CK N$11338 VDD p L=2u W=6u
        MN757 N$11338 N$11339 N$11099 GND n L=2u W=6u
        MN756 N$11333 CK GND GND n L=2u W=5u
        MP756 N$11333 CK VDD VDD p L=2u W=5u
        MN765 N$11339 CK GND GND n L=2u W=5u
        MN755 N$11337 N$11336 GND GND n L=2u W=6u
        MP755 N$11337 N$11336 VDD VDD p L=2u W=6u
        MN754 N$382 N$11337 GND GND n L=2u W=6u
        MP738 N$11328 N$11329 VDD VDD p L=2u W=6u
        MN724 N$11319 N$11318 GND GND n L=2u W=6u
        MN14 N$23 N$17 GND GND n L=2u W=6u
        MP313 N$346 N$344 VDD VDD p L=2u W=6u
        MN312 N$345 N$346 GND GND n L=2u W=6u
        MP312 N$345 N$346 VDD VDD p L=2u W=6u
        MN123 N$138 N$136 GND GND n L=2u W=3u
        MP127 N$136 GND N$135 VDD p L=2u W=3u
        MP126 N$136 N$120 N$132 VDD p L=2u W=3u
        MP125 N$135 N$388 N$132 VDD p L=2u W=3u
        MP124 N$132 N$388 VDD VDD p L=2u W=3u
        MN315 OUT8 N$11347 GND GND n L=2u W=5u
        MP315 GND N$348 OUT8 VDD p L=2u W=5u
        MP295 N$332 N$330 VDD VDD p L=2u W=6u
        MP349 N$14090 N$11347 N$397 VDD p L=2u W=5u
        MP348 N$331 N$14095 N$412 VDD p L=2u W=5u
        MN347 N$412 N$14095 N$14089 GND n L=2u W=5u
        MP347 N$14089 N$11347 N$412 VDD p L=2u W=5u
        MN346 N$376 N$11347 N$324 GND n L=2u W=5u
        MP346 N$324 N$14095 N$376 VDD p L=2u W=5u
        MN414 N$1661 N$11809 GND GND n L=2u W=3u
        MN413 N$1661 N$1673 GND GND n L=2u W=3u
        MN412 N$1661 N$1654 GND GND n L=2u W=3u
        MP422 N$1652 N$1653 N$1655 VDD p L=2u W=3u
        MP421 N$1655 N$1653 VDD VDD p L=2u W=3u
        MP420 N$1655 N$11561 VDD VDD p L=2u W=3u
        MP444 N$1628 N$1636 N$1629 VDD p L=2u W=3u
        MP443 N$1629 N$11786 N$1630 VDD p L=2u W=3u
        MN419 N$13038 N$1662 GND GND n L=2u W=3u
        MP419 N$13038 N$1662 VDD VDD p L=2u W=3u
        MN418 N$1662 N$11809 N$1660 GND n L=2u W=3u
        MN422 N$1651 N$1668 N$1649 GND n L=2u W=3u
        MN421 N$1649 N$11561 GND GND n L=2u W=3u
        MN420 N$1650 N$1651 GND GND n L=2u W=3u
        MP424 N$1651 N$11561 N$1652 VDD p L=2u W=3u
        MP423 N$1651 N$1668 N$1655 VDD p L=2u W=3u
        MP428 N$1647 N$1653 VDD VDD p L=2u W=3u
        MP427 N$1647 N$11561 VDD VDD p L=2u W=3u
        MN15 N$20 N$16 N$24 GND n L=2u W=6u
        MP538 N$1544 CK VDD VDD p L=2u W=5u
        MP765 N$11339 CK VDD VDD p L=2u W=5u
        MN764 N$11343 N$11342 GND GND n L=2u W=6u
        MP764 N$11343 N$11342 VDD VDD p L=2u W=6u
        MN763 N$11344 N$11343 GND GND n L=2u W=6u
        MP763 N$11344 N$11343 VDD VDD p L=2u W=6u
        MP762 N$11342 CK N$11344 VDD p L=2u W=6u
        MN762 N$11344 N$11339 N$11342 GND n L=2u W=6u
        MP761 N$11340 N$11339 N$11342 VDD p L=2u W=6u
        MN761 N$11342 CK N$11340 GND n L=2u W=6u
        MN760 N$11340 N$11341 GND GND n L=2u W=6u
        MP760 N$11340 N$11341 VDD VDD p L=2u W=6u
        MN539 N$1539 N$13857 GND GND n L=2u W=6u
        MP539 N$1539 N$13857 VDD VDD p L=2u W=6u
        MN538 N$1544 CK GND GND n L=2u W=5u
        MN537 N$11083 N$1540 GND GND n L=2u W=6u
        MP558 N$1521 CK N$1523 VDD p L=2u W=6u
        MN558 N$1523 N$1522 N$1521 GND n L=2u W=6u
        MN557 N$1525 N$1530 GND GND n L=2u W=5u
        MP563 N$1517 CK SK0 VDD p L=2u W=6u
        MP536 N$1554 N$11083 VDD VDD p L=2u W=6u
        MP535 N$1540 CK N$1554 VDD p L=2u W=6u
        MP770 N$11810 N$11802 VDD VDD p L=2u W=3u
        MN770 N$11810 N$11802 GND GND n L=2u W=3u
        MN520 N$1553 N$1558 GND GND n L=2u W=5u
        MN519 N$13857 N$1554 N$1553 GND n L=2u W=5u
        MP520 N$13857 N$1558 VDD VDD p L=2u W=5u
        MP519 N$13857 N$1554 VDD VDD p L=2u W=5u
        MP724 N$11319 N$11318 VDD VDD p L=2u W=6u
        MN723 N$14096 N$11319 GND GND n L=2u W=6u
        MN746 N$11345 N$11099 GND GND n L=2u W=5u
        MN745 N$11345 N$14096 GND GND n L=2u W=5u
        MN744 N$11345 N$382 GND GND n L=2u W=5u
        MP766 N$11345 N$11088 N$11108 VDD p L=2u W=5u
        MN522 N$1549 CK N$1552 GND n L=2u W=6u
        MP521 N$13650 CK N$1552 VDD p L=2u W=6u
        MP413 N$1665 N$1654 VDD VDD p L=2u W=3u
        MP412 N$1665 N$11809 VDD VDD p L=2u W=3u
        MN417 N$1662 N$1671 N$1661 GND n L=2u W=3u
        MN416 N$1659 N$1673 GND GND n L=2u W=3u
        MN415 N$1660 N$1654 N$1659 GND n L=2u W=3u
        MN499 N$1573 N$1572 N$1595 GND n L=2u W=6u
        MP504 N$1569 CK N$12429 VDD p L=2u W=6u
        MN504 N$12429 N$1572 N$1569 GND n L=2u W=6u
        MP472 N$13243 N$13447 VDD VDD p L=2u W=5u
        MN471 N$1595 N$13243 N$11786 GND n L=2u W=5u
        MP389 N$11780 CK VDD VDD p L=2u W=5u
        MP477 N$11561 N$13243 N$11816 VDD p L=2u W=5u
        MN476 N$11817 N$13243 N$11561 GND n L=2u W=5u
        MP476 N$11561 N$13447 N$11817 VDD p L=2u W=5u
        MN475 N$11817 N$13447 N$11786 GND n L=2u W=5u
        MP475 N$11786 N$13243 N$11817 VDD p L=2u W=5u
        MN389 N$11780 CK GND GND n L=2u W=5u
        MP480 N$1674 N$13447 N$1593 VDD p L=2u W=5u
        MN479 N$1593 N$13447 N$1654 GND n L=2u W=5u
        MP479 N$1654 N$13243 N$1593 VDD p L=2u W=5u
        MN478 N$11816 N$13243 N$1654 GND n L=2u W=5u
        MP478 N$1654 N$13447 N$11816 VDD p L=2u W=5u
        MN477 N$11816 N$13447 N$11561 GND n L=2u W=5u
        MP483 N$1584 N$1589 VDD VDD p L=2u W=6u
        MN518 N$1557 N$11083 GND GND n L=2u W=5u
        MN517 N$1557 N$1558 GND GND n L=2u W=5u
        MP524 N$1549 N$1548 VDD VDD p L=2u W=6u
        MN523 N$1548 N$1552 GND GND n L=2u W=6u
        MP523 N$1548 N$1552 VDD VDD p L=2u W=6u
        MP522 N$1552 N$1551 N$1549 VDD p L=2u W=6u
        MN500 N$1571 CK N$1573 GND n L=2u W=6u
        MN486 N$11571 N$1588 N$1583 GND n L=2u W=6u
        MP485 N$1585 N$1588 N$1583 VDD p L=2u W=6u
        MP469 N$13650 N$12835 N$1602 VDD p L=2u W=6u
        MN483 N$1584 N$1589 GND GND n L=2u W=6u
        MN461 N$13039 N$1611 GND GND n L=2u W=3u
        MP461 N$13039 N$1611 VDD VDD p L=2u W=3u
        MN473 N$13650 N$13039 GND GND n L=2u W=5u
        MP433 N$13037 N$1644 VDD VDD p L=2u W=3u
        MN432 N$1644 N$1668 N$1642 GND n L=2u W=3u
        MN431 N$1644 N$1651 N$1643 GND n L=2u W=3u
        MN430 N$1641 N$1653 GND GND n L=2u W=3u
        MN429 N$1642 N$11561 N$1641 GND n L=2u W=3u
        MN434 N$1633 N$1634 GND GND n L=2u W=3u
        MP438 N$1634 N$11786 N$1635 VDD p L=2u W=3u
        MP437 N$1634 N$1650 N$1638 VDD p L=2u W=3u
        MP436 N$1635 N$1636 N$1638 VDD p L=2u W=3u
        MP435 N$1638 N$1636 VDD VDD p L=2u W=3u
        MP434 N$1638 N$11786 VDD VDD p L=2u W=3u
        MP439 N$1633 N$1634 VDD VDD p L=2u W=3u
        MN439 N$1634 N$11786 N$1631 GND n L=2u W=3u
        MN438 N$1632 N$1636 GND GND n L=2u W=3u
        MN437 N$1631 N$1636 GND GND n L=2u W=3u
        MN436 N$1634 N$1650 N$1632 GND n L=2u W=3u
        MN470 N$1595 N$13447 N$1599 GND n L=2u W=5u
        MP470 N$1599 N$13243 N$1595 VDD p L=2u W=5u
        MN469 N$13650 N$12835 GND GND n L=2u W=6u
        MN468 N$13650 N$13037 GND GND n L=2u W=6u
        MN467 N$13650 N$13038 GND GND n L=2u W=6u
        MN541 N$1674 N$11813 N$1539 GND n L=2u W=5u
        MN472 N$13243 N$13447 GND GND n L=2u W=5u
        MN445 N$1627 N$1634 N$1626 GND n L=2u W=3u
        MN444 N$1624 N$1636 GND GND n L=2u W=3u
        MN443 N$1625 N$11786 N$1624 GND n L=2u W=3u
        MN388 N$11775 N$11777 GND GND n L=2u W=6u
        MP499 N$1595 CK N$1573 VDD p L=2u W=6u
        MP456 N$1614 N$1620 VDD VDD p L=2u W=3u
        MP455 N$1614 N$1599 VDD VDD p L=2u W=3u
        MP454 N$1614 N$1633 VDD VDD p L=2u W=3u
        MP453 N$13447 N$9715 VDD VDD p L=2u W=3u
        MN453 N$9715 N$1599 N$1615 GND n L=2u W=3u
        MN457 N$1609 N$1599 N$1608 GND n L=2u W=3u
        MN456 N$1610 N$1633 GND GND n L=2u W=3u
        MN440 N$1626 N$11786 GND GND n L=2u W=3u
        MN441 N$1626 N$1636 GND GND n L=2u W=3u
        MN442 N$1626 N$1650 GND GND n L=2u W=3u
        MN521 N$1552 N$1551 N$13650 GND n L=2u W=6u
        MP488 N$1581 N$1583 VDD VDD p L=2u W=6u
        MN487 N$11571 N$1581 GND GND n L=2u W=6u
        MP487 N$11571 N$1581 VDD VDD p L=2u W=6u
        MN507 N$1572 CK GND GND n L=2u W=5u
        MP507 N$1572 CK VDD VDD p L=2u W=5u
        MN506 N$12633 N$1569 GND GND n L=2u W=6u
        MP506 N$12633 N$1569 VDD VDD p L=2u W=6u
        MN435 N$1632 N$11786 GND GND n L=2u W=3u
        MP446 N$1627 N$1634 N$1630 VDD p L=2u W=3u
        MP445 N$1627 N$1650 N$1628 VDD p L=2u W=3u
        MN433 N$13037 N$1644 GND GND n L=2u W=3u
        MP429 N$1646 N$11561 N$1647 VDD p L=2u W=3u
        MP430 N$1645 N$1653 N$1646 VDD p L=2u W=3u
        MP591 SK3 N$1491 VDD VDD p L=2u W=6u
        MP590 N$1493 CK SK3 VDD p L=2u W=6u
        MN590 SK3 N$1497 N$1493 GND n L=2u W=6u
        MP589 N$1495 N$1497 N$1493 VDD p L=2u W=6u
        MN563 SK0 N$1522 N$1517 GND n L=2u W=6u
        MP562 N$1519 N$1522 N$1517 VDD p L=2u W=6u
        MN562 N$1517 CK N$1519 GND n L=2u W=6u
        MN155 N$174 N$390 GND GND n L=2u W=3u
        MN154 N$175 N$390 GND GND n L=2u W=3u
        MN198 N$222 N$14081 N$226 GND n L=2u W=3u
        MN197 N$225 N$395 GND GND n L=2u W=3u
        MN196 N$226 N$395 GND GND n L=2u W=3u
        MN195 N$222 N$207 N$225 GND n L=2u W=3u
        MN194 N$225 N$14081 GND GND n L=2u W=3u
        MP153 N$170 N$390 N$168 VDD p L=2u W=3u
        MP152 N$168 N$390 VDD VDD p L=2u W=3u
        MN94 N$94 N$90 GND GND n L=2u W=3u
        MP94 N$94 N$90 VDD VDD p L=2u W=3u
        MN93 N$90 GND N$92 GND n L=2u W=3u
        MN92 N$90 N$81 N$91 GND n L=2u W=3u
        MN91 N$93 N$385 GND GND n L=2u W=3u
        MN90 N$92 GND N$93 GND n L=2u W=3u
        MN89 N$91 GND GND GND n L=2u W=3u
        MP291 N$328 N$329 VDD VDD p L=2u W=6u
        MN290 N$329 N$326 GND GND n L=2u W=6u
        MP344 N$317 N$14095 N$411 VDD p L=2u W=5u
        MP289 N$326 N$327 N$328 VDD p L=2u W=6u
        MN289 N$328 CK N$326 GND n L=2u W=6u
        MP288 N$258 CK N$326 VDD p L=2u W=6u
        MP298 N$333 N$334 N$335 VDD p L=2u W=6u
        MN298 N$335 CK N$333 GND n L=2u W=6u
        MP87 N$87 GND VDD VDD p L=2u W=3u
        MP86 N$84 N$81 VDD VDD p L=2u W=3u
        MN86 N$81 GND N$86 GND n L=2u W=3u
        MN85 N$85 N$385 GND GND n L=2u W=3u
        MN113 N$121 N$387 GND GND n L=2u W=3u
        MN142 N$154 GND N$158 GND n L=2u W=3u
        MN141 N$157 N$389 GND GND n L=2u W=3u
        MN409 N$1666 N$1673 GND GND n L=2u W=3u
        MN408 N$1671 N$11809 N$1667 GND n L=2u W=3u
        MN455 N$1610 N$1620 GND GND n L=2u W=3u
        MN454 N$1610 N$1599 GND GND n L=2u W=3u
        MP460 N$1611 N$9715 N$1614 VDD p L=2u W=3u
        MP459 N$1611 N$1633 N$1612 VDD p L=2u W=3u
        MP458 N$1612 N$1620 N$1613 VDD p L=2u W=3u
        MN426 N$1643 N$11561 GND GND n L=2u W=3u
        MP432 N$1644 N$1651 N$1647 VDD p L=2u W=3u
        MP431 N$1644 N$1668 N$1645 VDD p L=2u W=3u
        MN266 N$310 N$306 N$309 GND n L=2u W=6u
        MP265 N$307 N$306 N$309 VDD p L=2u W=6u
        MN265 N$309 CK N$307 GND n L=2u W=6u
        MN264 N$307 N$308 GND GND n L=2u W=6u
        MP264 N$307 N$308 VDD VDD p L=2u W=6u
        MN263 N$308 N$305 GND GND n L=2u W=6u
        MP263 N$308 N$305 VDD VDD p L=2u W=6u
        MN240 N$417 N$420 GND GND n L=2u W=6u
        MP240 N$417 N$420 VDD VDD p L=2u W=6u
        MN205 N$230 N$207 N$232 GND n L=2u W=3u
        MN239 N$420 N$279 GND GND n L=2u W=6u
        MN238 N$420 N$386 GND GND n L=2u W=6u
        MP239 N$420 N$386 N$278 VDD p L=2u W=6u
        MP238 N$278 N$279 VDD VDD p L=2u W=6u
        MN258 N$384 N$304 GND GND n L=2u W=6u
        MP258 N$384 N$304 VDD VDD p L=2u W=6u
        MP257 N$302 CK N$384 VDD p L=2u W=6u
        MN257 N$384 N$299 N$302 GND n L=2u W=6u
        MN282 N$321 N$322 GND GND n L=2u W=6u
        MP282 N$321 N$322 VDD VDD p L=2u W=6u
        MN281 N$322 N$319 GND GND n L=2u W=6u
        MP501 N$1570 N$1573 VDD VDD p L=2u W=6u
        MP500 N$1573 N$1572 N$1571 VDD p L=2u W=6u
        MN532 N$1541 N$1545 GND GND n L=2u W=6u
        MP532 N$1541 N$1545 VDD VDD p L=2u W=6u
        MP531 N$1545 N$1544 N$1542 VDD p L=2u W=6u
        MN531 N$1542 CK N$1545 GND n L=2u W=6u
        MN536 N$1554 N$11083 GND GND n L=2u W=6u
        MP503 N$1571 N$1572 N$1569 VDD p L=2u W=6u
        MN503 N$1569 CK N$1571 GND n L=2u W=6u
        MN502 N$1571 N$1570 GND GND n L=2u W=6u
        MP276 N$317 N$318 VDD VDD p L=2u W=6u
        MP275 N$316 CK N$317 VDD p L=2u W=6u
        MN275 N$317 N$313 N$316 GND n L=2u W=6u
        MP274 N$314 N$313 N$316 VDD p L=2u W=6u
        MN274 N$316 CK N$314 GND n L=2u W=6u
        MN273 N$314 N$315 GND GND n L=2u W=6u
        MP273 N$314 N$315 VDD VDD p L=2u W=6u
        MN246 N$293 N$294 GND GND n L=2u W=6u
        MP246 N$293 N$294 VDD VDD p L=2u W=6u
        MP217 N$183 N$14095 N$250 VDD p L=2u W=5u
        MP245 N$294 N$291 VDD VDD p L=2u W=6u
        MP244 N$291 N$292 N$293 VDD p L=2u W=6u
        MN244 N$293 CK N$291 GND n L=2u W=6u
        MP243 N$237 CK N$291 VDD p L=2u W=6u
        MN243 N$291 N$292 N$237 GND n L=2u W=6u
        MP406 N$1675 N$1654 VDD VDD p L=2u W=3u
        MP262 N$305 N$306 N$307 VDD p L=2u W=6u
        MN262 N$307 CK N$305 GND n L=2u W=6u
        MP261 N$246 CK N$305 VDD p L=2u W=6u
        MP411 N$1668 N$1671 VDD VDD p L=2u W=3u
        MN411 N$1671 N$1654 N$1666 GND n L=2u W=3u
        MN410 N$1667 N$1673 GND GND n L=2u W=3u
        MN576 N$1506 N$1505 N$1504 GND n L=2u W=6u
        MN575 N$1513 CK GND GND n L=2u W=5u
        MP602 GND N$1557 N$1484 VDD p L=2u W=5u
        MN601 N$1484 N$1557 N$12429 GND n L=2u W=5u
        MN606 N$1475 N$1481 GND GND n L=2u W=3u
        MN605 N$1479 C N$1476 GND n L=2u W=3u
        MN604 N$1476 B0 GND GND n L=2u W=3u
        MN573 SK1 N$1507 GND GND n L=2u W=6u
        MP579 N$1503 N$1502 VDD VDD p L=2u W=6u
        MN578 N$1502 N$1506 GND GND n L=2u W=6u
        MP486 N$1583 CK N$11571 VDD p L=2u W=6u
        MN492 N$1577 N$1580 GND GND n L=2u W=6u
        MP492 N$1577 N$1580 VDD VDD p L=2u W=6u
        MP491 N$1580 N$1579 N$1578 VDD p L=2u W=6u
        MN491 N$1578 CK N$1580 GND n L=2u W=6u
        MP490 N$11816 CK N$1580 VDD p L=2u W=6u
        MN490 N$1580 N$1579 N$11816 GND n L=2u W=6u
        MN489 N$1588 CK GND GND n L=2u W=5u
        MP495 N$1576 CK N$11572 VDD p L=2u W=6u
        MN261 N$305 N$306 N$246 GND n L=2u W=6u
        MN260 N$299 CK GND GND n L=2u W=5u
        MP260 N$299 CK VDD VDD p L=2u W=5u
        MN259 N$304 N$302 GND GND n L=2u W=6u
        MP259 N$304 N$302 VDD VDD p L=2u W=6u
        MP498 N$1579 CK VDD VDD p L=2u W=5u
        MN497 N$1574 N$1576 GND GND n L=2u W=6u
        MP497 N$1574 N$1576 VDD VDD p L=2u W=6u
        MN496 N$11572 N$1574 GND GND n L=2u W=6u
        MP496 N$11572 N$1574 VDD VDD p L=2u W=6u
        MN501 N$1570 N$1573 GND GND n L=2u W=6u
        MN586 N$1495 CK N$1498 GND n L=2u W=6u
        MP585 N$1496 CK N$1498 VDD p L=2u W=6u
        MP618 N$1466 N$1465 VDD VDD p L=2u W=3u
        MP617 N$1466 B1 VDD VDD p L=2u W=3u
        MP623 N$1459 N$1477 VDD VDD p L=2u W=3u
        MP622 N$1462 N$1463 VDD VDD p L=2u W=3u
        MN622 N$1463 B1 N$1460 GND n L=2u W=3u
        MN589 N$1493 CK N$1495 GND n L=2u W=6u
        MN594 N$1488 N$1557 N$11571 GND n L=2u W=5u
        MP594 N$11571 N$1489 N$1488 VDD p L=2u W=5u
        MN561 N$1519 N$1518 GND GND n L=2u W=6u
        MP561 N$1519 N$1518 VDD VDD p L=2u W=6u
        MN566 N$1522 CK GND GND n L=2u W=5u
        MP566 N$1522 CK VDD VDD p L=2u W=5u
        MN565 N$1515 N$1517 GND GND n L=2u W=6u
        MP565 N$1515 N$1517 VDD VDD p L=2u W=6u
        MN564 SK0 N$1515 GND GND n L=2u W=6u
        MP564 SK0 N$1515 VDD VDD p L=2u W=6u
        MN245 N$294 N$291 GND GND n L=2u W=6u
        MN406 N$1668 N$1671 GND GND n L=2u W=3u
        MP410 N$1671 N$1654 N$1672 VDD p L=2u W=3u
        MP409 N$1671 N$11809 N$1675 VDD p L=2u W=3u
        MP408 N$1672 N$1673 N$1675 VDD p L=2u W=3u
        MP407 N$1675 N$1673 VDD VDD p L=2u W=3u
        MN567 N$1514 N$1513 N$1512 GND n L=2u W=6u
        MP573 SK1 N$1507 VDD VDD p L=2u W=6u
        MP572 N$1509 CK SK1 VDD p L=2u W=6u
        MN572 SK1 N$1513 N$1509 GND n L=2u W=6u
        MP571 N$1511 N$1513 N$1509 VDD p L=2u W=6u
        MN571 N$1509 CK N$1511 GND n L=2u W=6u
        MN570 N$1511 N$1510 GND GND n L=2u W=6u
        MN602 N$1484 N$1489 GND GND n L=2u W=5u
        MP635 N$1448 B2 N$1449 VDD p L=2u W=3u
        MP641 N$1442 N$1450 N$1443 VDD p L=2u W=3u
        MP640 N$1443 B2 N$1444 VDD p L=2u W=3u
        MP639 N$1444 N$1450 VDD VDD p L=2u W=3u
        MP638 N$1444 B2 VDD VDD p L=2u W=3u
        MN603 N$1477 N$1479 GND GND n L=2u W=3u
        MP607 N$1479 B0 N$1480 VDD p L=2u W=3u
        MP606 N$1479 C N$1482 VDD p L=2u W=3u
        MP578 N$1502 N$1506 VDD VDD p L=2u W=6u
        MP577 N$1506 N$1505 N$1503 VDD p L=2u W=6u
        MN577 N$1503 CK N$1506 GND n L=2u W=6u
        MP576 N$1504 CK N$1506 VDD p L=2u W=6u
        MP582 SK2 N$1499 VDD VDD p L=2u W=6u
        MP581 N$1501 CK SK2 VDD p L=2u W=6u
        MN581 SK2 N$1505 N$1501 GND n L=2u W=6u
        MP580 N$1503 N$1505 N$1501 VDD p L=2u W=6u
        MN580 N$1501 CK N$1503 GND n L=2u W=6u
        MN495 N$11572 N$1579 N$1576 GND n L=2u W=6u
        MP494 N$1578 N$1579 N$1576 VDD p L=2u W=6u
        MN494 N$1576 CK N$1578 GND n L=2u W=6u
        MN493 N$1578 N$1577 GND GND n L=2u W=6u
        MP493 N$1578 N$1577 VDD VDD p L=2u W=6u
        MN498 N$1579 CK GND GND n L=2u W=5u
        MP583 N$1499 N$1501 VDD VDD p L=2u W=6u
        MN582 SK2 N$1499 GND GND n L=2u W=6u
        MN588 N$1495 N$1494 GND GND n L=2u W=6u
        MP588 N$1495 N$1494 VDD VDD p L=2u W=6u
        MN587 N$1494 N$1498 GND GND n L=2u W=6u
        MP587 N$1494 N$1498 VDD VDD p L=2u W=6u
        MP586 N$1498 N$1497 N$1495 VDD p L=2u W=6u
        MP620 N$1463 N$1477 N$1466 VDD p L=2u W=3u
        MP619 N$1464 N$1465 N$1466 VDD p L=2u W=3u
        MN649 N$1431 N$1435 GND GND n L=2u W=3u
        MN648 N$1430 N$1435 GND GND n L=2u W=3u
        MN652 N$1425 N$1435 GND GND n L=2u W=3u
        MN651 N$1425 B3 GND GND n L=2u W=3u
        MP657 N$1426 N$1433 N$1429 VDD p L=2u W=3u
        MN621 N$1461 N$1465 GND GND n L=2u W=3u
        MN620 N$1460 N$1465 GND GND n L=2u W=3u
        MN619 N$1463 N$1477 N$1461 GND n L=2u W=3u
        MN593 N$1497 CK GND GND n L=2u W=5u
        MP593 N$1497 CK VDD VDD p L=2u W=5u
        MN592 N$1491 N$1493 GND GND n L=2u W=6u
        MP592 N$1491 N$1493 VDD VDD p L=2u W=6u
        MN597 N$1486 N$1557 N$11572 GND n L=2u W=5u
        MP597 N$11572 N$1489 N$1486 VDD p L=2u W=5u
        MN596 N$1489 N$1557 GND GND n L=2u W=5u
        MP570 N$1511 N$1510 VDD VDD p L=2u W=6u
        MN569 N$1510 N$1514 GND GND n L=2u W=6u
        MP569 N$1510 N$1514 VDD VDD p L=2u W=6u
        MP568 N$1514 N$1513 N$1511 VDD p L=2u W=6u
        MN568 N$1511 CK N$1514 GND n L=2u W=6u
        MP567 N$1512 CK N$1514 VDD p L=2u W=6u
        MN599 N$1485 N$1557 N$12632 GND n L=2u W=5u
        MP599 N$12632 N$1489 N$1485 VDD p L=2u W=5u
        MN598 N$1486 N$1489 GND GND n L=2u W=5u
        MP598 GND N$1557 N$1486 VDD p L=2u W=5u
        MP605 N$1480 N$1481 N$1482 VDD p L=2u W=3u
        MP604 N$1482 N$1481 VDD VDD p L=2u W=3u
        MP603 N$1482 B0 VDD VDD p L=2u W=3u
        MN632 N$1446 B2 GND GND n L=2u W=3u
        MN631 N$1447 N$1448 GND GND n L=2u W=3u
        MN667 N$1512 N$1416 N$1527 GND n L=2u W=5u
        MP667 N$1527 N$1557 N$1512 VDD p L=2u W=5u
        MN666 N$1512 N$1557 N$1486 GND n L=2u W=5u
        MP672 N$1467 N$1413 N$14097 VDD p L=2u W=5u
        MN671 N$1496 N$1416 N$1525 GND n L=2u W=5u
        MP637 N$1444 N$1462 VDD VDD p L=2u W=3u
        MP636 N$1447 N$1448 VDD VDD p L=2u W=3u
        MN636 N$1448 B2 N$1445 GND n L=2u W=3u
        MP611 N$1474 N$1481 VDD VDD p L=2u W=3u
        MP610 N$1474 B0 VDD VDD p L=2u W=3u
        MP609 N$1474 C VDD VDD p L=2u W=3u
        MP608 N$1477 N$1479 VDD VDD p L=2u W=3u
        MN608 N$1479 B0 N$1475 GND n L=2u W=3u
        MN607 N$1476 N$1481 GND GND n L=2u W=3u
        MN611 N$1470 C GND GND n L=2u W=3u
        MN610 N$1470 N$1481 GND GND n L=2u W=3u
        MN609 N$1470 B0 GND GND n L=2u W=3u
        MN579 N$1503 N$1502 GND GND n L=2u W=6u
        MN585 N$1498 N$1497 N$1496 GND n L=2u W=6u
        MN584 N$1505 CK GND GND n L=2u W=5u
        MP584 N$1505 CK VDD VDD p L=2u W=5u
        MN583 N$1499 N$1501 GND GND n L=2u W=6u
        MN615 N$1471 C N$1469 GND n L=2u W=3u
        MN614 N$1471 N$1479 N$1470 GND n L=2u W=3u
        MN613 N$1468 N$1481 GND GND n L=2u W=3u
        MN612 N$1469 B0 N$1468 GND n L=2u W=3u
        MN618 N$1461 B1 GND GND n L=2u W=3u
        MN617 N$1462 N$1463 GND GND n L=2u W=3u
        MP621 N$1463 B1 N$1464 VDD p L=2u W=3u
        MP650 COUTHK-SK N$1433 VDD VDD p L=2u W=3u
        MN650 N$1433 B3 N$1430 GND n L=2u W=3u
        MP684 N$1404 N$1403 VDD VDD p L=2u W=6u
        MN683 N$1403 N$1406 GND GND n L=2u W=6u
        MP683 N$1403 N$1406 VDD VDD p L=2u W=6u
        MP682 N$1406 N$14098 N$1404 VDD p L=2u W=6u
        MN682 N$1404 CK N$1406 GND n L=2u W=6u
        MP656 N$1426 N$1447 N$1427 VDD p L=2u W=3u
        MP655 N$1427 N$1435 N$1428 VDD p L=2u W=3u
        MP654 N$1428 B3 N$1429 VDD p L=2u W=3u
        MP629 N$1456 N$1463 N$1459 VDD p L=2u W=3u
        MP628 N$1456 N$1477 N$1457 VDD p L=2u W=3u
        MP627 N$1457 N$1465 N$1458 VDD p L=2u W=3u
        MP626 N$1458 B1 N$1459 VDD p L=2u W=3u
        MP625 N$1459 N$1465 VDD VDD p L=2u W=3u
        MP624 N$1459 B1 VDD VDD p L=2u W=3u
        MN629 N$1456 N$1477 N$1454 GND n L=2u W=3u
        MN628 N$1456 N$1463 N$1455 GND n L=2u W=3u
        MN627 N$1453 N$1465 GND GND n L=2u W=3u
        MP596 N$1489 N$1557 VDD VDD p L=2u W=5u
        MN595 N$1488 N$1489 GND GND n L=2u W=5u
        MP595 GND N$1557 N$1488 VDD p L=2u W=5u
        MP601 N$12429 N$1489 N$1484 VDD p L=2u W=5u
        MN600 N$1485 N$1489 GND GND n L=2u W=5u
        MP600 GND N$1557 N$1485 VDD p L=2u W=5u
        MP632 N$1451 N$1450 VDD VDD p L=2u W=3u
        MP631 N$1451 B2 VDD VDD p L=2u W=3u
        MN630 N$1452 N$1456 GND GND n L=2u W=3u
        MP630 N$1452 N$1456 VDD VDD p L=2u W=3u
        MN634 N$1445 N$1450 GND GND n L=2u W=3u
        MN633 N$1448 N$1462 N$1446 GND n L=2u W=3u
        MN668 N$1504 N$1557 N$1485 GND n L=2u W=5u
        MP668 N$1485 N$1416 N$1504 VDD p L=2u W=5u
        MN700 N$1392 CK N$1394 GND n L=2u W=6u
        MP699 N$1409 CK N$1394 VDD p L=2u W=6u
        MN699 N$1394 N$1393 N$1409 GND n L=2u W=6u
        MN698 N$1399 CK GND GND n L=2u W=5u
        MP698 N$1399 CK VDD VDD p L=2u W=5u
        MP671 N$1525 N$1557 N$1496 VDD p L=2u W=5u
        MN670 N$1496 N$1557 N$1484 GND n L=2u W=5u
        MN635 N$1446 N$1450 GND GND n L=2u W=3u
        MN640 N$1439 B2 N$1438 GND n L=2u W=3u
        MN639 N$1440 N$1462 GND GND n L=2u W=3u
        MN638 N$1440 N$1450 GND GND n L=2u W=3u
        MN637 N$1440 B2 GND GND n L=2u W=3u
        MP643 N$1441 N$1448 N$1444 VDD p L=2u W=3u
        MP642 N$1441 N$1462 N$1442 VDD p L=2u W=3u
        MP645 N$1436 B3 VDD VDD p L=2u W=3u
        MN644 N$1437 N$1441 GND GND n L=2u W=3u
        MP615 N$1471 N$1479 N$1474 VDD p L=2u W=3u
        MP614 N$1471 C N$1472 VDD p L=2u W=3u
        MP613 N$1472 N$1481 N$1473 VDD p L=2u W=3u
        MP612 N$1473 B0 N$1474 VDD p L=2u W=3u
        MN616 N$1467 N$1471 GND GND n L=2u W=3u
        MP616 N$1467 N$1471 VDD VDD p L=2u W=3u
        MN645 COUTHK-SK N$1433 GND GND n L=2u W=3u
        MP649 N$1433 B3 N$1434 VDD p L=2u W=3u
        MP648 N$1433 N$1447 N$1436 VDD p L=2u W=3u
        MP647 N$1434 N$1435 N$1436 VDD p L=2u W=3u
        MP646 N$1436 N$1435 VDD VDD p L=2u W=3u
        MP652 N$1429 B3 VDD VDD p L=2u W=3u
        MP651 N$1429 N$1447 VDD VDD p L=2u W=3u
        MP679 N$1422 N$1413 N$1408 VDD p L=2u W=5u
        MN684 N$1404 N$1403 GND GND n L=2u W=6u
        MP716 N$1387 CK VDD VDD p L=2u W=5u
        MN715 N$1383 N$1384 GND GND n L=2u W=6u
        MP715 N$1383 N$1384 VDD VDD p L=2u W=6u
        MN714 N$14092 N$1383 GND GND n L=2u W=6u
        MP714 N$14092 N$1383 VDD VDD p L=2u W=6u
        MP688 N$1401 N$1402 VDD VDD p L=2u W=6u
        MN687 N$14046 N$1401 GND GND n L=2u W=6u
        MP687 N$14046 N$1401 VDD VDD p L=2u W=6u
        MP653 N$1429 N$1435 VDD VDD p L=2u W=3u
        MP658 N$1422 N$1426 VDD VDD p L=2u W=3u
        MN657 N$1426 N$1447 N$1424 GND n L=2u W=3u
        MN656 N$1426 N$1433 N$1425 GND n L=2u W=3u
        MN655 N$1423 N$1435 GND GND n L=2u W=3u
        MN654 N$1424 B3 N$1423 GND n L=2u W=3u
        MN653 N$1425 N$1447 GND GND n L=2u W=3u
        MP661 N$1435 N$1484 VDD VDD p L=2u W=3u
        MN660 N$1465 N$1486 GND GND n L=2u W=3u
        MN626 N$1454 B1 N$1453 GND n L=2u W=3u
        MN625 N$1455 N$1477 GND GND n L=2u W=3u
        MN624 N$1455 N$1465 GND GND n L=2u W=3u
        MN623 N$1455 B1 GND GND n L=2u W=3u
        MP634 N$1448 N$1462 N$1451 VDD p L=2u W=3u
        MP633 N$1449 N$1450 N$1451 VDD p L=2u W=3u
        MN665 N$1416 N$1557 GND GND n L=2u W=5u
        MP665 N$1416 N$1557 VDD VDD p L=2u W=5u
        MN664 N$1521 N$1416 N$1529 GND n L=2u W=5u
        MP664 N$1529 N$1557 N$1521 VDD p L=2u W=5u
        MN663 N$1521 N$1557 N$1488 GND n L=2u W=5u
        MP669 N$1526 N$1557 N$1504 VDD p L=2u W=5u
        MP556 N$12632 N$1530 N$1525 VDD p L=2u W=5u
        MN555 N$1526 N$1530 GND GND n L=2u W=5u
        MP555 GND N$1539 N$1526 VDD p L=2u W=5u
        MN554 N$1526 N$1539 N$11572 GND n L=2u W=5u
        MN560 N$1518 N$1523 GND GND n L=2u W=6u
        MP560 N$1518 N$1523 VDD VDD p L=2u W=6u
        MP559 N$1523 N$1522 N$1519 VDD p L=2u W=6u
        MN559 N$1519 CK N$1523 GND n L=2u W=6u
        MP489 N$1588 CK VDD VDD p L=2u W=5u
        MN488 N$1581 N$1583 GND GND n L=2u W=6u
        MN340 N$410 N$11347 N$384 GND n L=2u W=5u
        MP340 N$384 N$14095 N$410 VDD p L=2u W=5u
        MN339 N$410 N$14095 N$14085 GND n L=2u W=5u
        MP339 N$14085 N$11347 N$410 VDD p L=2u W=5u
        MP358 P2 N$409 N$387 VDD p L=2u W=5u
        MN358 N$387 N$14096 P2 GND n L=2u W=5u
        MP355 N$409 N$14096 VDD VDD p L=2u W=5u
        MN355 N$409 N$14096 GND GND n L=2u W=5u
        MN678 N$1409 N$1413 GND GND n L=2u W=5u
        MP678 GND N$1557 N$1409 VDD p L=2u W=5u
        MN677 N$1409 N$1557 N$1437 GND n L=2u W=5u
        MP677 N$1437 N$1413 N$1409 VDD p L=2u W=5u
        MN676 N$1410 N$1413 GND GND n L=2u W=5u
        MP676 GND N$1557 N$1410 VDD p L=2u W=5u
        MN708 N$1388 N$1387 N$1408 GND n L=2u W=6u
        MN707 N$1393 CK GND GND n L=2u W=5u
        MN713 N$14092 N$1387 N$1384 GND n L=2u W=6u
        MP712 N$1386 N$1387 N$1384 VDD p L=2u W=6u
        MN712 N$1384 CK N$1386 GND n L=2u W=6u
        MN711 N$1386 N$1385 GND GND n L=2u W=6u
        MP711 N$1386 N$1385 VDD VDD p L=2u W=6u
        MN511 N$13874 N$13996 GND GND n L=2u W=3u
        MN510 N$13875 N$13996 GND GND n L=2u W=3u
        MN509 N$13870 GND N$13874 GND n L=2u W=3u
        MN508 N$13874 N$14084 GND GND n L=2u W=3u
        MN474 N$13873 N$13870 GND GND n L=2u W=3u
        MP511 N$13870 N$14084 N$13869 VDD p L=2u W=3u
        MP510 N$13870 GND N$13868 VDD p L=2u W=3u
        MP509 N$13869 N$13996 N$13868 VDD p L=2u W=3u
        MP508 N$13868 N$13996 VDD VDD p L=2u W=3u
        MP474 N$13868 N$14084 VDD VDD p L=2u W=3u
        MP400 N$11799 N$11794 VDD VDD p L=2u W=3u
        MP399 N$11799 N$1674 VDD VDD p L=2u W=3u
        MP398 N$11799 C VDD VDD p L=2u W=3u
        MP397 N$11809 N$11796 VDD VDD p L=2u W=3u
        MN397 N$11796 N$1674 N$11798 GND n L=2u W=3u
        MN396 N$11797 N$11794 GND GND n L=2u W=3u
        MN395 N$11798 N$11794 GND GND n L=2u W=3u
        MN394 N$11796 C N$11797 GND n L=2u W=3u
        MN393 N$11797 N$1674 GND GND n L=2u W=3u
        MN235 N$421 N$275 GND GND n L=2u W=6u
        MN234 N$421 N$385 GND GND n L=2u W=6u
        MP235 N$421 N$385 N$274 VDD p L=2u W=6u
        MP234 N$274 N$275 VDD VDD p L=2u W=6u
        MP553 GND N$1539 N$1527 VDD p L=2u W=5u
        MN552 N$1527 N$1539 N$11571 GND n L=2u W=5u
        MP552 N$11571 N$1530 N$1527 VDD p L=2u W=5u
        MN551 N$1530 N$1539 GND GND n L=2u W=5u
        MP557 GND N$1539 N$1525 VDD p L=2u W=5u
        MN556 N$1525 N$1539 N$12632 GND n L=2u W=5u
        MP783 N$13889 N$13887 VDD VDD p L=2u W=3u
        MN783 N$13887 N$14085 N$13891 GND n L=2u W=3u
        MN782 N$13890 N$14000 GND GND n L=2u W=3u
        MN781 N$13891 N$14000 GND GND n L=2u W=3u
        MN780 N$13887 N$13873 N$13890 GND n L=2u W=3u
        MN779 N$13890 N$14085 GND GND n L=2u W=3u
        MN778 N$13889 N$13887 GND GND n L=2u W=3u
        MP782 N$13887 N$14085 N$13886 VDD p L=2u W=3u
        MP781 N$13887 N$13873 N$13885 VDD p L=2u W=3u
        MP780 N$13886 N$14000 N$13885 VDD p L=2u W=3u
        MP779 N$13885 N$14000 VDD VDD p L=2u W=3u
        MP778 N$13885 N$14085 VDD VDD p L=2u W=3u
        MN777 OUT0 N$13879 GND GND n L=2u W=3u
        MP777 OUT0 N$13879 VDD VDD p L=2u W=3u
        MN776 N$13879 GND N$13881 GND n L=2u W=3u
        MN775 N$13879 N$13870 N$13880 GND n L=2u W=3u
        MN774 N$13882 N$13996 GND GND n L=2u W=3u
        MN574 N$1507 N$1509 GND GND n L=2u W=6u
        MP575 N$1513 CK VDD VDD p L=2u W=5u
        MP554 N$11572 N$1530 N$1526 VDD p L=2u W=5u
        MN553 N$1527 N$1530 GND GND n L=2u W=5u
        MP774 N$13878 N$13996 N$13877 VDD p L=2u W=3u
        MP516 N$13877 N$14084 N$13876 VDD p L=2u W=3u
        MP515 N$13876 N$13996 VDD VDD p L=2u W=3u
        MP514 N$13876 N$14084 VDD VDD p L=2u W=3u
        MP513 N$13876 GND VDD VDD p L=2u W=3u
        MP512 N$13873 N$13870 VDD VDD p L=2u W=3u
        MN512 N$13870 N$14084 N$13875 GND n L=2u W=3u
        MP799 N$13908 N$14086 VDD VDD p L=2u W=3u
        MP798 N$13908 N$13889 VDD VDD p L=2u W=3u
        MP797 N$13905 N$13903 VDD VDD p L=2u W=3u
        MN797 N$13903 N$14086 N$13907 GND n L=2u W=3u
        MN796 N$13906 N$14001 GND GND n L=2u W=3u
        MN795 N$13907 N$14001 GND GND n L=2u W=3u
        MN794 N$13903 N$13889 N$13906 GND n L=2u W=3u
        MN793 N$13906 N$14086 GND GND n L=2u W=3u
        MN792 N$13905 N$13903 GND GND n L=2u W=3u
        MP796 N$13903 N$14086 N$13902 VDD p L=2u W=3u
        MP795 N$13903 N$13889 N$13901 VDD p L=2u W=3u
        MP794 N$13902 N$14001 N$13901 VDD p L=2u W=3u
        MP793 N$13901 N$14001 VDD VDD p L=2u W=3u
        MP792 N$13901 N$14086 VDD VDD p L=2u W=3u
        MN791 OUT1 N$13895 GND GND n L=2u W=3u
        MP791 OUT1 N$13895 VDD VDD p L=2u W=3u
        MN790 N$13895 N$13873 N$13897 GND n L=2u W=3u
        MN392 N$11809 N$11796 GND GND n L=2u W=3u
        MP396 N$11796 N$1674 N$11795 VDD p L=2u W=3u
        MP395 N$11796 C N$11793 VDD p L=2u W=3u
        MP394 N$11795 N$11794 N$11793 VDD p L=2u W=3u
        MP393 N$11793 N$11794 VDD VDD p L=2u W=3u
        MP392 N$11793 N$1674 VDD VDD p L=2u W=3u
        MP790 N$13895 N$13887 N$13892 VDD p L=2u W=3u
        MP789 N$13895 N$13873 N$13894 VDD p L=2u W=3u
        MP788 N$13894 N$14000 N$13893 VDD p L=2u W=3u
        MP787 N$13893 N$14085 N$13892 VDD p L=2u W=3u
        MP786 N$13892 N$14000 VDD VDD p L=2u W=3u
        MP785 N$13892 N$14085 VDD VDD p L=2u W=3u
        MP784 N$13892 N$13873 VDD VDD p L=2u W=3u
        MP815 N$13925 N$14087 N$13924 VDD p L=2u W=3u
        MP814 N$13924 N$14002 VDD VDD p L=2u W=3u
        MP813 N$13924 N$14087 VDD VDD p L=2u W=3u
        MP812 N$13924 N$13905 VDD VDD p L=2u W=3u
        MP811 N$13921 N$13919 VDD VDD p L=2u W=3u
        MN811 N$13919 N$14087 N$13923 GND n L=2u W=3u
        MN810 N$13922 N$14002 GND GND n L=2u W=3u
        MN809 N$13923 N$14002 GND GND n L=2u W=3u
        MN808 N$13919 N$13905 N$13922 GND n L=2u W=3u
        MN807 N$13922 N$14087 GND GND n L=2u W=3u
        MN806 N$13921 N$13919 GND GND n L=2u W=3u
        MP810 N$13919 N$14087 N$13918 VDD p L=2u W=3u
        MP809 N$13919 N$13905 N$13917 VDD p L=2u W=3u
        MP808 N$13918 N$14002 N$13917 VDD p L=2u W=3u
        MP807 N$13917 N$14002 VDD VDD p L=2u W=3u
        MP806 N$13917 N$14087 VDD VDD p L=2u W=3u
        MN805 OUT2 N$13911 GND GND n L=2u W=3u
        MN516 N$13881 N$14084 N$13882 GND n L=2u W=3u
        MN515 N$13880 GND GND GND n L=2u W=3u
        MN514 N$13880 N$13996 GND GND n L=2u W=3u
        MN513 N$13880 N$14084 GND GND n L=2u W=3u
        MP776 N$13879 N$13870 N$13876 VDD p L=2u W=3u
        MP775 N$13879 GND N$13878 VDD p L=2u W=3u
        MN799 N$13912 N$14001 GND GND n L=2u W=3u
        MN798 N$13912 N$14086 GND GND n L=2u W=3u
        MP804 N$13911 N$13903 N$13908 VDD p L=2u W=3u
        MP803 N$13911 N$13889 N$13910 VDD p L=2u W=3u
        MP802 N$13910 N$14001 N$13909 VDD p L=2u W=3u
        MP801 N$13909 N$14086 N$13908 VDD p L=2u W=3u
        MP800 N$13908 N$14001 VDD VDD p L=2u W=3u
        MP831 N$13943 N$13921 N$13942 VDD p L=2u W=3u
        MP830 N$13942 N$14003 N$13941 VDD p L=2u W=3u
        MP829 N$13941 N$14088 N$13940 VDD p L=2u W=3u
        MP828 N$13940 N$14003 VDD VDD p L=2u W=3u
        MP827 N$13940 N$14088 VDD VDD p L=2u W=3u
        MP826 N$13940 N$13921 VDD VDD p L=2u W=3u
        MP825 N$13937 N$13935 VDD VDD p L=2u W=3u
        MN825 N$13935 N$14088 N$13939 GND n L=2u W=3u
        MN824 N$13938 N$14003 GND GND n L=2u W=3u
        MN823 N$13939 N$14003 GND GND n L=2u W=3u
        MN822 N$13935 N$13921 N$13938 GND n L=2u W=3u
        MN821 N$13938 N$14088 GND GND n L=2u W=3u
        MN820 N$13937 N$13935 GND GND n L=2u W=3u
        MP824 N$13935 N$14088 N$13934 VDD p L=2u W=3u
        MP823 N$13935 N$13921 N$13933 VDD p L=2u W=3u
        MP822 N$13934 N$14003 N$13933 VDD p L=2u W=3u
        MP821 N$13933 N$14003 VDD VDD p L=2u W=3u
        MP820 N$13933 N$14088 VDD VDD p L=2u W=3u
        MN789 N$13895 N$13887 N$13896 GND n L=2u W=3u
        MN788 N$13898 N$14000 GND GND n L=2u W=3u
        MN787 N$13897 N$14085 N$13898 GND n L=2u W=3u
        MN786 N$13896 N$13873 GND GND n L=2u W=3u
        MN785 N$13896 N$14000 GND GND n L=2u W=3u
        MN784 N$13896 N$14085 GND GND n L=2u W=3u
        MN815 N$13929 N$14087 N$13930 GND n L=2u W=3u
        MN814 N$13928 N$13905 GND GND n L=2u W=3u
        MN813 N$13928 N$14002 GND GND n L=2u W=3u
        MN812 N$13928 N$14087 GND GND n L=2u W=3u
        MP818 N$13927 N$13919 N$13924 VDD p L=2u W=3u
        MP817 N$13927 N$13905 N$13926 VDD p L=2u W=3u
        MP816 N$13926 N$14002 N$13925 VDD p L=2u W=3u
        MN840 N$13960 N$14089 GND GND n L=2u W=3u
        MP846 N$13959 N$13951 N$13956 VDD p L=2u W=3u
        MP845 N$13959 N$13937 N$13958 VDD p L=2u W=3u
        MP844 N$13958 N$14004 N$13957 VDD p L=2u W=3u
        MP843 N$13957 N$14089 N$13956 VDD p L=2u W=3u
        MP842 N$13956 N$14004 VDD VDD p L=2u W=3u
        MP841 N$13956 N$14089 VDD VDD p L=2u W=3u
        MP840 N$13956 N$13937 VDD VDD p L=2u W=3u
        MP839 N$13953 N$13951 VDD VDD p L=2u W=3u
        MN839 N$13951 N$14089 N$13955 GND n L=2u W=3u
        MN838 N$13954 N$14004 GND GND n L=2u W=3u
        MN837 N$13955 N$14004 GND GND n L=2u W=3u
        MN836 N$13951 N$13937 N$13954 GND n L=2u W=3u
        MN835 N$13954 N$14089 GND GND n L=2u W=3u
        MN834 N$13953 N$13951 GND GND n L=2u W=3u
        MP838 N$13951 N$14089 N$13950 VDD p L=2u W=3u
        MP837 N$13951 N$13937 N$13949 VDD p L=2u W=3u
        MP836 N$13950 N$14004 N$13949 VDD p L=2u W=3u
        MP835 N$13949 N$14004 VDD VDD p L=2u W=3u
        MP805 OUT2 N$13911 VDD VDD p L=2u W=3u
        MN804 N$13911 N$13889 N$13913 GND n L=2u W=3u
        MN803 N$13911 N$13903 N$13912 GND n L=2u W=3u
        MN802 N$13914 N$14001 GND GND n L=2u W=3u
        MN801 N$13913 N$14086 N$13914 GND n L=2u W=3u
        MN800 N$13912 N$13889 GND GND n L=2u W=3u
        MN831 N$13943 N$13935 N$13944 GND n L=2u W=3u
        MN830 N$13946 N$14003 GND GND n L=2u W=3u
        MN829 N$13945 N$14088 N$13946 GND n L=2u W=3u
        MN828 N$13944 N$13921 GND GND n L=2u W=3u
        MN827 N$13944 N$14003 GND GND n L=2u W=3u
        MN826 N$13944 N$14088 GND GND n L=2u W=3u
        MP832 N$13943 N$13935 N$13940 VDD p L=2u W=3u
        MN856 N$13976 N$13953 GND GND n L=2u W=3u
        MN855 N$13976 N$14005 GND GND n L=2u W=3u
        MN854 N$13976 N$14090 GND GND n L=2u W=3u
        MP860 N$13975 N$13967 N$13972 VDD p L=2u W=3u
        MP859 N$13975 N$13953 N$13974 VDD p L=2u W=3u
        MP858 N$13974 N$14005 N$13973 VDD p L=2u W=3u
        MP857 N$13973 N$14090 N$13972 VDD p L=2u W=3u
        MP856 N$13972 N$14005 VDD VDD p L=2u W=3u
        MP855 N$13972 N$14090 VDD VDD p L=2u W=3u
        MP854 N$13972 N$13953 VDD VDD p L=2u W=3u
        MP853 N$13969 N$13967 VDD VDD p L=2u W=3u
        MN853 N$13967 N$14090 N$13971 GND n L=2u W=3u
        MN852 N$13970 N$14005 GND GND n L=2u W=3u
        MN851 N$13971 N$14005 GND GND n L=2u W=3u
        MN850 N$13967 N$13953 N$13970 GND n L=2u W=3u
        MN849 N$13970 N$14090 GND GND n L=2u W=3u
        MN848 N$13969 N$13967 GND GND n L=2u W=3u
        MP852 N$13967 N$14090 N$13966 VDD p L=2u W=3u
        MP851 N$13967 N$13953 N$13965 VDD p L=2u W=3u
        MN819 OUT3 N$13927 GND GND n L=2u W=3u
        MP819 OUT3 N$13927 VDD VDD p L=2u W=3u
        MN818 N$13927 N$13905 N$13929 GND n L=2u W=3u
        MN817 N$13927 N$13919 N$13928 GND n L=2u W=3u
        MN816 N$13930 N$14002 GND GND n L=2u W=3u
        MP847 OUT5 N$13959 VDD VDD p L=2u W=3u
        MN846 N$13959 N$13937 N$13961 GND n L=2u W=3u
        MN845 N$13959 N$13951 N$13960 GND n L=2u W=3u
        MN844 N$13962 N$14004 GND GND n L=2u W=3u
        MN843 N$13961 N$14089 N$13962 GND n L=2u W=3u
        MN842 N$13960 N$13937 GND GND n L=2u W=3u
        MN841 N$13960 N$14004 GND GND n L=2u W=3u
        MN872 N$13994 N$14007 GND GND n L=2u W=3u
        MN871 N$13993 N$14091 N$13994 GND n L=2u W=3u
        MN870 N$13992 N$13969 GND GND n L=2u W=3u
        MN869 N$13992 N$14007 GND GND n L=2u W=3u
        MN868 N$13992 N$14091 GND GND n L=2u W=3u
        MP874 N$13991 N$13983 N$13988 VDD p L=2u W=3u
        MP873 N$13991 N$13969 N$13990 VDD p L=2u W=3u
        MP872 N$13990 N$14007 N$13989 VDD p L=2u W=3u
        MP871 N$13989 N$14091 N$13988 VDD p L=2u W=3u
        MP870 N$13988 N$14007 VDD VDD p L=2u W=3u
        MP869 N$13988 N$14091 VDD VDD p L=2u W=3u
        MP868 N$13988 N$13969 VDD VDD p L=2u W=3u
        MP867 CARRY_OUT N$13983 VDD VDD p L=2u W=3u
        MN867 N$13983 N$14091 N$13987 GND n L=2u W=3u
        MN866 N$13986 N$14007 GND GND n L=2u W=3u
        MN865 N$13987 N$14007 GND GND n L=2u W=3u
        MN864 N$13983 N$13969 N$13986 GND n L=2u W=3u
        MN863 N$13986 N$14091 GND GND n L=2u W=3u
        MN862 CARRY_OUT N$13983 GND GND n L=2u W=3u
        MP834 N$13949 N$14089 VDD VDD p L=2u W=3u
        MN833 OUT4 N$13943 GND GND n L=2u W=3u
        MP833 OUT4 N$13943 VDD VDD p L=2u W=3u
        MN832 N$13943 N$13921 N$13945 GND n L=2u W=3u
        MN861 OUT6 N$13975 GND GND n L=2u W=3u
        MP861 OUT6 N$13975 VDD VDD p L=2u W=3u
        MN860 N$13975 N$13953 N$13977 GND n L=2u W=3u
        MN859 N$13975 N$13967 N$13976 GND n L=2u W=3u
        MN858 N$13978 N$14005 GND GND n L=2u W=3u
        MN857 N$13977 N$14090 N$13978 GND n L=2u W=3u
        MP923 N$14018 SK2 N$14009 VDD p L=2u W=5u
        MN922 N$14010 SK2 N$14017 GND n L=2u W=5u
        MP922 N$14017 N$14015 N$14010 VDD p L=2u W=5u
        MP928 N$14012 N$14006 N$14007 VDD p L=2u W=5u
        MN927 N$14007 N$14006 N$14016 GND n L=2u W=5u
        MP927 N$14016 SK3 N$14007 VDD p L=2u W=5u
        MN926 N$14008 SK2 GND GND n L=2u W=5u
        MP926 GND N$14015 N$14008 VDD p L=2u W=5u
        MN925 N$14008 N$14015 N$14017 GND n L=2u W=5u
        MP925 N$14017 SK2 N$14008 VDD p L=2u W=5u
        MP931 N$14011 N$14006 N$14005 VDD p L=2u W=5u
        MN930 N$14005 N$14006 N$14014 GND n L=2u W=5u
        MP930 N$14014 SK3 N$14005 VDD p L=2u W=5u
        MN929 N$14006 SK3 GND GND n L=2u W=5u
        MP929 N$14006 SK3 VDD VDD p L=2u W=5u
        MN928 N$14007 SK3 N$14012 GND n L=2u W=5u
        MP934 N$14012 SK3 N$14003 VDD p L=2u W=5u
        MN933 N$14004 SK3 N$14010 GND n L=2u W=5u
        MP933 N$14010 N$14006 N$14004 VDD p L=2u W=5u
        MN900 N$14021 N$14024 N$14031 GND n L=2u W=5u
        MP900 N$14031 SK1 N$14021 VDD p L=2u W=5u
        MN899 N$14022 SK1 N$14031 GND n L=2u W=5u
        MN905 N$14019 SK1 N$14028 GND n L=2u W=5u
        MP905 N$14028 N$14024 N$14019 VDD p L=2u W=5u
        MN904 N$14019 N$14024 N$14029 GND n L=2u W=5u
        MP904 N$14029 SK1 N$14019 VDD p L=2u W=5u
        MN903 N$14020 SK1 N$14029 GND n L=2u W=5u
        MP903 N$14029 N$14024 N$14020 VDD p L=2u W=5u
        MN902 N$14020 N$14024 N$14030 GND n L=2u W=5u
        MN908 N$14017 N$14024 N$14027 GND n L=2u W=5u
        MP908 N$14027 SK1 N$14017 VDD p L=2u W=5u
        MN907 N$14018 SK1 N$14027 GND n L=2u W=5u
        MP939 GND N$14006 N$14001 VDD p L=2u W=5u
        MN938 N$14001 N$14006 N$14010 GND n L=2u W=5u
        MP938 N$14010 SK3 N$14001 VDD p L=2u W=5u
        MP944 N$11083 N$13857 N$14040 VDD p L=2u W=5u
        MN943 N$13996 SK3 GND GND n L=2u W=5u
        MP943 GND N$14006 N$13996 VDD p L=2u W=5u
        MN942 N$13996 N$14006 N$14008 GND n L=2u W=5u
        MP942 N$14008 SK3 N$13996 VDD p L=2u W=5u
        MN941 N$14000 SK3 GND GND n L=2u W=5u
        MP941 GND N$14006 N$14000 VDD p L=2u W=5u
        MN946 N$13997 N$11083 GND GND n L=2u W=5u
        MP947 N$13997 N$11347 N$13998 VDD p L=2u W=5u
        MP946 N$13998 N$11083 VDD VDD p L=2u W=5u
        MN945 N$14040 N$13857 N$13999 GND n L=2u W=5u
        MP945 N$13999 N$1539 N$14040 VDD p L=2u W=5u
        MN944 N$14040 N$1539 N$11083 GND n L=2u W=5u
        MN948 N$13999 N$13997 GND GND n L=2u W=5u
        MP948 N$13999 N$13997 VDD VDD p L=2u W=5u
        MN947 N$13997 N$11347 GND GND n L=2u W=5u
        MN916 N$14013 SK2 N$14020 GND n L=2u W=5u
        MP916 N$14020 N$14015 N$14013 VDD p L=2u W=5u
        MN915 N$14013 N$14015 N$14022 GND n L=2u W=5u
        MN921 N$14010 N$14015 N$14019 GND n L=2u W=5u
        MP921 N$14019 SK2 N$14010 VDD p L=2u W=5u
        MN920 N$14011 SK2 N$14018 GND n L=2u W=5u
        MP920 N$14018 N$14015 N$14011 VDD p L=2u W=5u
        MN919 N$14011 N$14015 N$14020 GND n L=2u W=5u
        MP919 N$14020 SK2 N$14011 VDD p L=2u W=5u
        MN918 N$14012 SK2 N$14019 GND n L=2u W=5u
        MN924 N$14009 SK2 GND GND n L=2u W=5u
        MP924 GND N$14015 N$14009 VDD p L=2u W=5u
        MN923 N$14009 N$14015 N$14018 GND n L=2u W=5u
        MP130 N$141 GND VDD VDD p L=2u W=3u
        MP129 N$141 N$120 VDD VDD p L=2u W=3u
        MP128 N$138 N$136 VDD VDD p L=2u W=3u
        MP172 N$193 N$14079 VDD VDD p L=2u W=3u
        MP201 N$227 N$395 VDD VDD p L=2u W=3u
        MP200 N$227 N$14081 VDD VDD p L=2u W=3u
        MP199 N$227 N$207 VDD VDD p L=2u W=3u
        MP198 COUT N$222 VDD VDD p L=2u W=3u
        MN223 N$258 N$265 N$217 GND n L=2u W=5u
        MP223 N$217 N$14095 N$258 VDD p L=2u W=5u
        MN222 N$258 N$14095 N$200 GND n L=2u W=5u
        MP222 N$200 N$265 N$258 VDD p L=2u W=5u
        MP418 N$1662 N$1671 N$1665 VDD p L=2u W=3u
        MP417 N$1662 N$11809 N$1663 VDD p L=2u W=3u
        MP416 N$1663 N$1673 N$1664 VDD p L=2u W=3u
        MP415 N$1664 N$1654 N$1665 VDD p L=2u W=3u
        MN299 N$336 N$333 GND GND n L=2u W=6u
        MP299 N$336 N$333 VDD VDD p L=2u W=6u
        MP266 N$309 CK N$310 VDD p L=2u W=6u
        MP232 N$112 N$14095 N$271 VDD p L=2u W=5u
        MN231 N$271 N$14095 N$94 GND n L=2u W=5u
        MP231 N$94 N$265 N$271 VDD p L=2u W=5u
        MN407 N$1667 N$1654 GND GND n L=2u W=3u
        MP302 N$337 CK N$338 VDD p L=2u W=6u
        MP303 N$338 N$339 VDD VDD p L=2u W=6u
        MN206 N$1179 N$230 GND GND n L=2u W=3u
        MP206 N$1179 N$230 VDD VDD p L=2u W=3u
        MN145 N$163 N$138 GND GND n L=2u W=3u
        MN204 N$230 N$222 N$231 GND n L=2u W=3u
        MN203 N$233 N$395 GND GND n L=2u W=3u
        MN202 N$232 N$14081 N$233 GND n L=2u W=3u
        MN201 N$231 N$207 GND GND n L=2u W=3u
        MN200 N$231 N$395 GND GND n L=2u W=3u
        MN237 N$275 N$386 GND GND n L=2u W=6u
        MP237 N$275 N$386 VDD VDD p L=2u W=6u
        MN236 N$419 N$421 GND GND n L=2u W=6u
        MP236 N$419 N$421 VDD VDD p L=2u W=6u
        MP256 N$300 N$299 N$302 VDD p L=2u W=6u
        MN288 N$326 N$327 N$258 GND n L=2u W=6u
        MN287 N$320 CK GND GND n L=2u W=5u
        MN193 COUT N$222 GND GND n L=2u W=3u
        MP197 N$222 N$14081 N$221 VDD p L=2u W=3u
        MP151 N$168 N$14078 VDD VDD p L=2u W=3u
        MP131 N$141 N$388 VDD VDD p L=2u W=3u
        MN122 N$130 N$126 GND GND n L=2u W=3u
        MP122 N$130 N$126 VDD VDD p L=2u W=3u
        MN121 N$126 N$102 N$128 GND n L=2u W=3u
        MN120 N$126 N$118 N$127 GND n L=2u W=3u
        MN119 N$129 N$387 GND GND n L=2u W=3u
        MN118 N$128 GND N$129 GND n L=2u W=3u
        MN88 N$91 N$385 GND GND n L=2u W=3u
        MN87 N$91 GND GND GND n L=2u W=3u
        MP93 N$90 N$81 N$87 VDD p L=2u W=3u
        MP121 N$126 N$118 N$123 VDD p L=2u W=3u
        MP120 N$126 N$102 N$125 VDD p L=2u W=3u
        MP119 N$125 N$387 N$124 VDD p L=2u W=3u
        MP118 N$124 GND N$123 VDD p L=2u W=3u
        MP117 N$123 N$387 VDD VDD p L=2u W=3u
        MN546 N$11561 N$11813 N$11572 GND n L=2u W=5u
        MP546 N$11572 RST N$11561 VDD p L=2u W=5u
        MN545 N$11561 RST GND GND n L=2u W=5u
        MP545 GND N$11813 N$11561 VDD p L=2u W=5u
        MN544 N$1654 N$11813 N$11571 GND n L=2u W=5u
        MP544 N$11571 RST N$1654 VDD p L=2u W=5u
        MN543 N$1654 RST GND GND n L=2u W=5u
        MN542 N$11813 RST GND GND n L=2u W=5u
        MP543 GND N$11813 N$1654 VDD p L=2u W=5u
        MP377 N$11790 CK N$1539 VDD p L=2u W=6u
        MN377 N$1539 N$11789 N$11790 GND n L=2u W=6u
        MN169 N$191 N$392 GND GND n L=2u W=3u
        MN211 N$242 N$265 N$148 GND n L=2u W=5u
        MP211 N$148 N$14095 N$242 VDD p L=2u W=5u
        MN210 N$242 N$14095 N$130 GND n L=2u W=5u
        MP210 N$130 N$265 N$242 VDD p L=2u W=5u
        MN170 N$188 N$14079 N$192 GND n L=2u W=3u
        MP168 N$188 N$173 N$185 VDD p L=2u W=3u
        MP167 N$187 N$392 N$185 VDD p L=2u W=3u
        MN108 N$112 N$108 GND GND n L=2u W=3u
        MP108 N$112 N$108 VDD VDD p L=2u W=3u
        MN107 N$108 N$84 N$110 GND n L=2u W=3u
        MN106 N$108 N$100 N$109 GND n L=2u W=3u
        MN105 N$111 N$386 GND GND n L=2u W=3u
        MN104 N$110 GND N$111 GND n L=2u W=3u
        MN103 N$109 N$84 GND GND n L=2u W=3u
        MP316 N$361 N$11347 OUT8 VDD p L=2u W=5u
        MP309 N$342 N$343 VDD VDD p L=2u W=6u
        MN330 N$14089 N$348 N$331 GND n L=2u W=5u
        MP308 N$343 N$340 VDD VDD p L=2u W=6u
        MP307 N$340 N$341 N$342 VDD p L=2u W=6u
        MN307 N$342 CK N$340 GND n L=2u W=6u
        MP306 N$266 CK N$340 VDD p L=2u W=6u
        MN306 N$340 N$341 N$266 GND n L=2u W=6u
        MP101 N$105 N$84 VDD VDD p L=2u W=3u
        MP100 N$102 N$100 VDD VDD p L=2u W=3u
        MN100 N$100 GND N$104 GND n L=2u W=3u
        MN99 N$103 N$386 GND GND n L=2u W=3u
        MN128 N$136 GND N$140 GND n L=2u W=3u
        MP156 N$173 N$171 VDD VDD p L=2u W=3u
        MN156 N$171 N$14078 N$175 GND n L=2u W=3u
        MP320 GND N$348 N$14085 VDD p L=2u W=5u
        MN329 N$14089 N$11347 GND GND n L=2u W=5u
        MP329 GND N$348 N$14089 VDD p L=2u W=5u
        MP185 N$210 N$190 VDD VDD p L=2u W=3u
        MP184 N$207 N$205 VDD VDD p L=2u W=3u
        MN184 N$205 N$14080 N$209 GND n L=2u W=3u
        MN183 N$208 N$394 GND GND n L=2u W=3u
        MN182 N$209 N$394 GND GND n L=2u W=3u
        MN181 N$205 N$190 N$208 GND n L=2u W=3u
        MN180 N$208 N$14080 GND GND n L=2u W=3u
        MN95 N$102 N$100 GND GND n L=2u W=3u
        MP99 N$100 GND N$99 VDD p L=2u W=3u
        MP12 N$15 N$17 VDD VDD p L=2u W=6u
        MN692 N$1397 N$1400 GND GND n L=2u W=6u
        MP692 N$1397 N$1400 VDD VDD p L=2u W=6u
        MP109 N$114 GND VDD VDD p L=2u W=3u
        MN233 N$265 N$14095 GND GND n L=2u W=5u
        MP233 N$265 N$14095 VDD VDD p L=2u W=5u
        MN189 N$216 N$394 GND GND n L=2u W=3u
        MP110 N$114 N$387 VDD VDD p L=2u W=3u
        MN208 N$237 N$265 N$130 GND n L=2u W=5u
        MP208 N$130 N$14095 N$237 VDD p L=2u W=5u
        MN207 N$237 N$14095 N$112 GND n L=2u W=5u
        MP375 N$11783 N$11782 VDD VDD p L=2u W=6u
        MN374 N$11782 N$11784 GND GND n L=2u W=6u
        MP374 N$11782 N$11784 VDD VDD p L=2u W=6u
        MP373 N$11784 N$11789 N$11783 VDD p L=2u W=6u
        MN373 N$11783 CK N$11784 GND n L=2u W=6u
        MP372 N$11570 CK N$11784 VDD p L=2u W=6u
        MP64 N$286 N$287 VDD VDD p L=2u W=6u
        MN63 N$287 N$282 GND GND n L=2u W=6u
        MP63 N$287 N$282 VDD VDD p L=2u W=6u
        MN64 N$286 N$287 GND GND n L=2u W=6u
        MN65 N$288 CK N$286 GND n L=2u W=6u
        MP181 N$204 N$394 N$202 VDD p L=2u W=3u
        MN136 N$148 N$144 GND GND n L=2u W=3u
        MP136 N$148 N$144 VDD VDD p L=2u W=3u
        MN135 N$144 N$120 N$146 GND n L=2u W=3u
        MN134 N$144 N$136 N$145 GND n L=2u W=3u
        MN133 N$147 N$388 GND GND n L=2u W=3u
        MN102 N$109 N$386 GND GND n L=2u W=3u
        MN101 N$109 GND GND GND n L=2u W=3u
        MP290 N$329 N$326 VDD VDD p L=2u W=6u
        MP92 N$90 GND N$89 VDD p L=2u W=3u
        MP91 N$89 N$385 N$88 VDD p L=2u W=3u
        MP90 N$88 GND N$87 VDD p L=2u W=3u
        MP89 N$87 N$385 VDD VDD p L=2u W=3u
        MP88 N$87 GND VDD VDD p L=2u W=3u
        MP116 N$123 GND VDD VDD p L=2u W=3u
        MP115 N$123 N$102 VDD VDD p L=2u W=3u
        MP114 N$120 N$118 VDD VDD p L=2u W=3u
        MN114 N$118 GND N$122 GND n L=2u W=3u
        MP142 N$156 N$154 VDD VDD p L=2u W=3u
        MP171 N$193 N$173 VDD VDD p L=2u W=3u
        MP170 N$190 N$188 VDD VDD p L=2u W=3u
        MN423 N$1648 N$1653 GND GND n L=2u W=3u
        MN428 N$1643 N$1668 GND GND n L=2u W=3u
        MN427 N$1643 N$1653 GND GND n L=2u W=3u
        MN277 N$318 N$316 GND GND n L=2u W=6u
        MP277 N$318 N$316 VDD VDD p L=2u W=6u
        MN276 N$317 N$318 GND GND n L=2u W=6u
        MP250 N$297 N$295 VDD VDD p L=2u W=6u
        MN249 N$296 N$297 GND GND n L=2u W=6u
        MP249 N$296 N$297 VDD VDD p L=2u W=6u
        MP248 N$295 CK N$296 VDD p L=2u W=6u
        MN248 N$296 N$292 N$295 GND n L=2u W=6u
        MP247 N$293 N$292 N$295 VDD p L=2u W=6u
        MN247 N$295 CK N$293 GND n L=2u W=6u
        MP280 N$319 N$320 N$321 VDD p L=2u W=6u
        MN217 N$250 N$265 N$183 GND n L=2u W=5u
        MN190 N$213 N$205 N$214 GND n L=2u W=3u
        MN216 N$250 N$14095 N$166 GND n L=2u W=5u
        MP216 N$166 N$265 N$250 VDD p L=2u W=5u
        MN425 N$1651 N$11561 N$1648 GND n L=2u W=3u
        MN424 N$1649 N$1653 GND GND n L=2u W=3u
        MP281 N$322 N$319 VDD VDD p L=2u W=6u
        MN242 N$283 CK GND GND n L=2u W=5u
        MP242 N$283 CK VDD VDD p L=2u W=5u
        MN68 N$290 N$288 GND GND n L=2u W=6u
        MP68 N$290 N$288 VDD VDD p L=2u W=6u
        MN272 N$315 N$312 GND GND n L=2u W=6u
        MP304 N$339 N$337 VDD VDD p L=2u W=6u
        MN303 N$338 N$339 GND GND n L=2u W=6u
        MN279 N$319 N$320 N$254 GND n L=2u W=6u
        MN278 N$313 CK GND GND n L=2u W=5u
        MP278 N$313 CK VDD VDD p L=2u W=5u
        MP283 N$321 N$320 N$323 VDD p L=2u W=6u
        MN283 N$323 CK N$321 GND n L=2u W=6u
        MN250 N$297 N$295 GND GND n L=2u W=6u
        MN220 N$254 N$265 N$200 GND n L=2u W=5u
        MP220 N$200 N$14095 N$254 VDD p L=2u W=5u
        MN219 N$254 N$14095 N$183 GND n L=2u W=5u
        MP219 N$183 N$265 N$254 VDD p L=2u W=5u
        MN280 N$321 CK N$319 GND n L=2u W=6u
        MP279 N$254 CK N$319 VDD p L=2u W=6u
        MN286 N$325 N$323 GND GND n L=2u W=6u
        MP192 N$217 N$213 VDD VDD p L=2u W=3u
        MN191 N$213 N$190 N$215 GND n L=2u W=3u
        MN130 N$145 N$388 GND GND n L=2u W=3u
        MN174 N$198 N$14079 N$199 GND n L=2u W=3u
        MN173 N$197 N$173 GND GND n L=2u W=3u
        MN172 N$197 N$392 GND GND n L=2u W=3u
        MN171 N$197 N$14079 GND GND n L=2u W=3u
        MP177 N$196 N$188 N$193 VDD p L=2u W=3u
        MP287 N$320 CK VDD VDD p L=2u W=5u
        MN214 N$246 N$265 N$166 GND n L=2u W=5u
        MP214 N$166 N$14095 N$246 VDD p L=2u W=5u
        MN213 N$246 N$14095 N$148 GND n L=2u W=5u
        MN256 N$302 CK N$300 GND n L=2u W=6u
        MN255 N$300 N$301 GND GND n L=2u W=6u
        MN139 N$154 N$138 N$157 GND n L=2u W=3u
        MN168 N$192 N$392 GND GND n L=2u W=3u
        MN167 N$188 N$173 N$191 GND n L=2u W=3u
        MN166 N$191 N$14079 GND GND n L=2u W=3u
        MN165 N$190 N$188 GND GND n L=2u W=3u
        MP169 N$188 N$14079 N$187 VDD p L=2u W=3u
        MP138 N$150 N$389 VDD VDD p L=2u W=3u
        MP137 N$150 GND VDD VDD p L=2u W=3u
        MP319 N$296 N$11347 N$14084 VDD p L=2u W=5u
        MN318 N$14084 N$11347 GND GND n L=2u W=5u
        MP318 GND N$348 N$14084 VDD p L=2u W=5u
        MN317 N$348 N$11347 GND GND n L=2u W=5u
        MP317 N$348 N$11347 VDD VDD p L=2u W=5u
        MN316 OUT8 N$348 N$361 GND n L=2u W=5u
        MN331 N$14090 N$11347 GND GND n L=2u W=5u
        MP331 GND N$348 N$14090 VDD p L=2u W=5u
        MN547 N$11786 RST GND GND n L=2u W=5u
        MP547 GND N$11813 N$11786 VDD p L=2u W=5u
        MN140 N$158 N$389 GND GND n L=2u W=3u
        MP527 N$1558 N$1546 VDD VDD p L=2u W=6u
        MN401 N$11804 N$1674 N$11805 GND n L=2u W=3u
        MN451 N$1615 N$1620 GND GND n L=2u W=3u
        MN450 N$9715 N$1633 N$1616 GND n L=2u W=3u
        MN449 N$1616 N$1599 GND GND n L=2u W=3u
        MN448 N$13447 N$9715 GND GND n L=2u W=3u
        MP452 N$9715 N$1599 N$1619 VDD p L=2u W=3u
        MP451 N$9715 N$1633 N$1622 VDD p L=2u W=3u
        MP457 N$1613 N$1599 N$1614 VDD p L=2u W=3u
        MN351 N$396 N$14095 N$14091 GND n L=2u W=5u
        MP351 N$14091 N$11347 N$396 VDD p L=2u W=5u
        MN731 N$11099 N$11321 N$11324 GND n L=2u W=6u
        MP731 N$11324 CK N$11099 VDD p L=2u W=6u
        MP732 N$11099 N$11325 VDD VDD p L=2u W=6u
        MP721 N$11316 N$11315 N$11318 VDD p L=2u W=6u
        MN721 N$11318 CK N$11316 GND n L=2u W=6u
        MN720 N$11316 N$11317 GND GND n L=2u W=6u
        MP720 N$11316 N$11317 VDD VDD p L=2u W=6u
        MN719 N$11317 N$11314 GND GND n L=2u W=6u
        MP719 N$11317 N$11314 VDD VDD p L=2u W=6u
        MP718 N$11314 N$11315 N$11316 VDD p L=2u W=6u
        MN718 N$11316 CK N$11314 GND n L=2u W=6u
        MP717 N$382 CK N$11314 VDD p L=2u W=6u
        MN752 N$11336 CK N$11334 GND n L=2u W=6u
        MP752 N$11334 N$11333 N$11336 VDD p L=2u W=6u
        MN753 N$382 N$11333 N$11336 GND n L=2u W=6u
        MN352 N$396 N$11347 N$345 GND n L=2u W=5u
        MP352 N$345 N$14095 N$396 VDD p L=2u W=5u
        MP83 N$80 N$385 N$77 VDD p L=2u W=3u
        MN226 N$262 N$265 N$1179 GND n L=2u W=5u
        MP226 N$1179 N$14095 N$262 VDD p L=2u W=5u
        MN225 N$262 N$14095 N$217 GND n L=2u W=5u
        MN67 N$361 N$290 GND GND n L=2u W=6u
        MP272 N$315 N$312 VDD VDD p L=2u W=6u
        MP163 N$179 N$171 N$176 VDD p L=2u W=3u
        MP162 N$179 N$156 N$178 VDD p L=2u W=3u
        MN526 N$1558 N$1551 N$1547 GND n L=2u W=6u
        MP525 N$1549 N$1551 N$1547 VDD p L=2u W=6u
        MN525 N$1547 CK N$1549 GND n L=2u W=6u
        MN524 N$1549 N$1548 GND GND n L=2u W=6u
        MP530 N$13447 CK N$1545 VDD p L=2u W=6u
        MN530 N$1545 N$1544 N$13447 GND n L=2u W=6u
        MN529 N$1551 CK GND GND n L=2u W=6u
        MP529 N$1551 CK VDD VDD p L=2u W=6u
        MN528 N$1546 N$1547 GND GND n L=2u W=6u
        MP528 N$1546 N$1547 VDD VDD p L=2u W=6u
        MN527 N$1558 N$1546 GND GND n L=2u W=6u
        MN533 N$1542 N$1541 GND GND n L=2u W=6u
        MP533 N$1542 N$1541 VDD VDD p L=2u W=6u
        MP473 N$13651 N$13039 VDD VDD p L=2u W=5u
        MN548 N$11786 N$11813 N$12632 GND n L=2u W=5u
        MP526 N$1547 CK N$1558 VDD p L=2u W=6u
        MP548 N$12632 RST N$11786 VDD p L=2u W=5u
        MP482 N$1589 N$1588 N$1585 VDD p L=2u W=6u
        MN482 N$1585 CK N$1589 GND n L=2u W=6u
        MP481 N$1593 CK N$1589 VDD p L=2u W=6u
        MN481 N$1589 N$1588 N$1593 GND n L=2u W=6u
        MN480 N$1593 N$13243 N$1674 GND n L=2u W=5u
        MN769 N$11802 C N$11804 GND n L=2u W=3u
        MN400 N$11803 C GND GND n L=2u W=3u
        MN399 N$11803 N$11794 GND GND n L=2u W=3u
        MN398 N$11803 N$1674 GND GND n L=2u W=3u
        MP769 N$11802 N$11796 N$11799 VDD p L=2u W=3u
        MP768 N$11802 C N$11801 VDD p L=2u W=3u
        MP402 N$11801 N$11794 N$11800 VDD p L=2u W=3u
        MP401 N$11800 N$1674 N$11799 VDD p L=2u W=3u
        MN459 N$1611 N$9715 N$1610 GND n L=2u W=3u
        MN458 N$1608 N$1620 GND GND n L=2u W=3u
        MN464 N$1620 GND GND GND n L=2u W=3u
        MP464 N$1620 GND VDD VDD p L=2u W=3u
        MN463 N$1653 B2 GND GND n L=2u W=3u
        MP463 N$1653 B2 VDD VDD p L=2u W=3u
        MN462 N$1673 B1 GND GND n L=2u W=3u
        MP462 N$1673 B1 VDD VDD p L=2u W=3u
        MN460 N$1611 N$1633 N$1609 GND n L=2u W=3u
        MN466 N$13650 N$11810 GND GND n L=2u W=6u
        MP484 N$1585 N$1584 VDD VDD p L=2u W=6u
        MP468 N$1602 N$13037 N$1603 VDD p L=2u W=6u
        MP467 N$1603 N$13038 N$1604 VDD p L=2u W=6u
        MP466 N$1604 N$11810 N$13651 VDD p L=2u W=6u
        MN465 N$1636 B3 GND GND n L=2u W=3u
        MP465 N$1636 B3 VDD VDD p L=2u W=3u
        MP471 N$11786 N$13447 N$1595 VDD p L=2u W=5u
        MP426 N$1647 N$1668 VDD VDD p L=2u W=3u
        MP425 N$1650 N$1651 VDD VDD p L=2u W=3u
        MP541 N$1539 RST N$1674 VDD p L=2u W=5u
        MN540 N$1674 RST A5 GND n L=2u W=5u
        MP540 A5 N$11813 N$1674 VDD p L=2u W=5u
        MP414 N$1665 N$1673 VDD VDD p L=2u W=3u
        MP442 N$1630 N$1636 VDD VDD p L=2u W=3u
        MP441 N$1630 N$11786 VDD VDD p L=2u W=3u
        MP440 N$1630 N$1650 VDD VDD p L=2u W=3u
        MP537 N$11083 N$1540 VDD VDD p L=2u W=6u
        MP534 N$1542 N$1544 N$1540 VDD p L=2u W=6u
        MN535 N$1554 N$1544 N$1540 GND n L=2u W=6u
        MN534 N$1540 CK N$1542 GND n L=2u W=6u
        MP888 GND N$14037 N$14029 VDD p L=2u W=5u
        MN887 N$14029 N$14037 P3 GND n L=2u W=5u
        MP896 N$14035 SK1 N$14023 VDD p L=2u W=5u
        MN895 N$14024 SK1 GND GND n L=2u W=5u
        MP895 N$14024 SK1 VDD VDD p L=2u W=5u
        MN894 N$14025 SK1 N$14035 GND n L=2u W=5u
        MP894 N$14035 N$14024 N$14025 VDD p L=2u W=5u
        MN893 N$14025 N$14024 N$14039 GND n L=2u W=5u
        MP899 N$14031 N$14024 N$14022 VDD p L=2u W=5u
        MN898 N$14022 N$14024 N$14033 GND n L=2u W=5u
        MP898 N$14033 SK1 N$14022 VDD p L=2u W=5u
        MN897 N$14023 SK1 N$14033 GND n L=2u W=5u
        MP897 N$14033 N$14024 N$14023 VDD p L=2u W=5u
        MN896 N$14023 N$14024 N$14035 GND n L=2u W=5u
        MP902 N$14030 SK1 N$14020 VDD p L=2u W=5u
        MN901 N$14021 SK1 N$14030 GND n L=2u W=5u
        MP901 N$14030 N$14024 N$14021 VDD p L=2u W=5u
        MP866 N$13983 N$14091 N$13982 VDD p L=2u W=3u
        MP865 N$13983 N$13969 N$13981 VDD p L=2u W=3u
        MP864 N$13982 N$14007 N$13981 VDD p L=2u W=3u
        MP863 N$13981 N$14007 VDD VDD p L=2u W=3u
        MP862 N$13981 N$14091 VDD VDD p L=2u W=3u
        MP878 N$14037 N$14040 VDD VDD p L=2u W=5u
        MN877 N$14039 N$14040 GND GND n L=2u W=5u
        MN888 N$14029 N$14040 GND GND n L=2u W=5u
        MP877 GND N$14037 N$14039 VDD p L=2u W=5u
        MN876 N$14039 N$14037 GND GND n L=2u W=5u
        MP876 GND N$14040 N$14039 VDD p L=2u W=5u
        MN906 N$14018 N$14024 N$14028 GND n L=2u W=5u
        MP906 N$14028 SK1 N$14018 VDD p L=2u W=5u
        MP912 N$14015 SK2 VDD VDD p L=2u W=5u
        MN911 N$14016 SK2 N$14022 GND n L=2u W=5u
        MP911 N$14022 N$14015 N$14016 VDD p L=2u W=5u
        MN910 N$14016 N$14015 N$14025 GND n L=2u W=5u
        MP910 N$14025 SK2 N$14016 VDD p L=2u W=5u
        MN909 N$14017 SK1 GND GND n L=2u W=5u
        MP909 GND N$14024 N$14017 VDD p L=2u W=5u
        MP915 N$14022 SK2 N$14013 VDD p L=2u W=5u
        MN914 N$14014 SK2 N$14021 GND n L=2u W=5u
        MP914 N$14021 N$14015 N$14014 VDD p L=2u W=5u
        MN913 N$14014 N$14015 N$14023 GND n L=2u W=5u
        MP913 N$14023 SK2 N$14014 VDD p L=2u W=5u
        MN912 N$14015 SK2 GND GND n L=2u W=5u
        MP918 N$14019 N$14015 N$14012 VDD p L=2u W=5u
        MN917 N$14012 N$14015 N$14021 GND n L=2u W=5u
        MP917 N$14021 SK2 N$14012 VDD p L=2u W=5u
        MP882 GND N$14037 N$14033 VDD p L=2u W=5u
        MN881 N$14033 N$14037 GND GND n L=2u W=5u
        MP881 GND N$14040 N$14033 VDD p L=2u W=5u
        MP887 P3 N$14040 N$14029 VDD p L=2u W=5u
        MN886 N$14030 N$14040 GND GND n L=2u W=5u
        MP886 GND N$14037 N$14030 VDD p L=2u W=5u
        MN885 N$14030 N$14037 P4 GND n L=2u W=5u
        MP885 P4 N$14040 N$14030 VDD p L=2u W=5u
        MN884 N$14031 N$14040 GND GND n L=2u W=5u
        MP907 N$14027 N$14024 N$14018 VDD p L=2u W=5u
        MP890 GND N$14037 N$14028 VDD p L=2u W=5u
        MN889 N$14028 N$14037 P2 GND n L=2u W=5u
        MP889 P2 N$14040 N$14028 VDD p L=2u W=5u
        MN376 N$11790 CK N$11783 GND n L=2u W=6u
        MN375 N$11783 N$11782 GND GND n L=2u W=6u
        MP381 N$11817 CK N$11781 VDD p L=2u W=6u
        MN381 N$11781 N$11780 N$11817 GND n L=2u W=6u
        MN380 N$11789 CK GND GND n L=2u W=5u
        MP380 N$11789 CK VDD VDD p L=2u W=5u
        MN379 N$11787 N$11790 GND GND n L=2u W=6u
        MP379 N$11787 N$11790 VDD VDD p L=2u W=6u
        MN384 N$11779 N$11778 GND GND n L=2u W=6u
        MP384 N$11779 N$11778 VDD VDD p L=2u W=6u
        MN383 N$11778 N$11781 GND GND n L=2u W=6u
        MP376 N$11783 N$11789 N$11790 VDD p L=2u W=6u
        MN892 N$14027 N$14040 GND GND n L=2u W=5u
        MP893 N$14039 SK1 N$14025 VDD p L=2u W=5u
        MP892 GND N$14037 N$14027 VDD p L=2u W=5u
        MN891 N$14027 N$14037 P1 GND n L=2u W=5u
        MN932 N$14004 N$14006 N$14013 GND n L=2u W=5u
        MP932 N$14013 SK3 N$14004 VDD p L=2u W=5u
        MN931 N$14005 SK3 N$14011 GND n L=2u W=5u
        MN937 N$14002 SK3 N$14008 GND n L=2u W=5u
        MP937 N$14008 N$14006 N$14002 VDD p L=2u W=5u
        MN936 N$14002 N$14006 N$14011 GND n L=2u W=5u
        MP936 N$14011 SK3 N$14002 VDD p L=2u W=5u
        MN935 N$14003 SK3 N$14009 GND n L=2u W=5u
        MP935 N$14009 N$14006 N$14003 VDD p L=2u W=5u
        MN934 N$14003 N$14006 N$14012 GND n L=2u W=5u
        MN940 N$14000 N$14006 N$14009 GND n L=2u W=5u
        MP940 N$14009 SK3 N$14000 VDD p L=2u W=5u
        MN939 N$14001 SK3 GND GND n L=2u W=5u
        MP743 N$11327 CK VDD VDD p L=2u W=5u
        MN741 N$11088 N$11331 GND GND n L=2u W=6u
        MN743 N$11327 CK GND GND n L=2u W=5u
        MN361 N$388 N$409 N$374 GND n L=2u W=5u
        MP753 N$11336 CK N$382 VDD p L=2u W=6u
        MN2 N$6 N$3 GND GND n L=2u W=6u
        MN1 N$2 ADD_ONE N$6 GND n L=2u W=6u
        MP2 N$2 ADD_ONE VDD VDD p L=2u W=6u
        MP1 N$2 N$3 VDD VDD p L=2u W=6u
        MP742 N$11331 N$11330 VDD VDD p L=2u W=6u
        MP754 N$382 N$11337 VDD VDD p L=2u W=6u
        MP241 N$279 N$385 VDD VDD p L=2u W=6u
        MP405 N$1180 N$1177 VDD VDD p L=2u W=5u
        MN241 N$279 N$385 GND GND n L=2u W=6u
        MN742 N$11331 N$11330 GND GND n L=2u W=6u
        MN405 N$1180 N$1177 GND GND n L=2u W=5u
        MP323 N$310 N$11347 N$14086 VDD p L=2u W=5u
        MP403 N$1176 N$1179 VDD VDD p L=2u W=5u
        MN323 N$14086 N$348 N$310 GND n L=2u W=5u
        MP404 N$1177 GND N$1176 VDD p L=2u W=5u
        MN325 N$14087 N$348 N$317 GND n L=2u W=5u
        MP19 N$25 N$20 VDD VDD p L=2u W=6u
        MN18 N$22 N$17 GND GND n L=2u W=6u
        MP18 N$22 N$17 VDD VDD p L=2u W=6u
        MN17 N$21 N$16 GND GND n L=2u W=6u
        MP17 N$21 N$16 VDD VDD p L=2u W=6u
        MN16 N$24 N$22 GND GND n L=2u W=6u
        MN21 N$27 N$14 N$29 GND n L=2u W=6u
        MP229 N$1180 N$14095 N$266 VDD p L=2u W=5u
        MN229 N$266 N$265 N$1180 GND n L=2u W=5u
        MN324 N$14087 N$11347 GND GND n L=2u W=5u
        MP357 N$372 N$14096 N$386 VDD p L=2u W=5u
        MN356 N$386 N$14096 P1 GND n L=2u W=5u
        MN6 N$12 N$10 GND GND n L=2u W=6u
        MN5 N$8 N$3 N$12 GND n L=2u W=6u
        MN4 N$11 ADD_ONE GND GND n L=2u W=6u
        MN3 N$8 N$9 N$11 GND n L=2u W=6u
        MN368 N$394 N$14096 GND GND n L=2u W=5u
        MP368 GND N$409 N$394 VDD p L=2u W=5u
        MN367 N$392 N$409 N$412 GND n L=2u W=5u
        MP367 N$412 N$14096 N$392 VDD p L=2u W=5u
        MN366 N$392 N$14096 GND GND n L=2u W=5u
        MP366 GND N$409 N$392 VDD p L=2u W=5u
        MP447 N$12835 N$1627 VDD VDD p L=2u W=3u
        MP449 N$1622 N$1620 VDD VDD p L=2u W=3u
        MP369 N$397 N$14096 N$394 VDD p L=2u W=5u
        MN452 N$1616 N$1620 GND GND n L=2u W=3u
        MN447 N$12835 N$1627 GND GND n L=2u W=3u
        MP448 N$1622 N$1599 VDD VDD p L=2u W=3u
        MN446 N$1627 N$1650 N$1625 GND n L=2u W=3u
        MN61 N$282 N$283 N$271 GND n L=2u W=6u
        MN228 N$266 N$14095 N$1179 GND n L=2u W=5u
        MP6 N$8 ADD_ONE N$7 VDD p L=2u W=6u
        MP96 N$96 N$386 VDD VDD p L=2u W=3u
        MP95 N$96 GND VDD VDD p L=2u W=3u
        MP228 N$1179 N$265 N$266 VDD p L=2u W=5u
        MP750 N$11335 N$11332 VDD VDD p L=2u W=6u
        MP10 N$14 N$2 VDD VDD p L=2u W=6u
        MN9 N$13 N$8 GND GND n L=2u W=6u
        MP9 N$13 N$8 VDD VDD p L=2u W=6u
        MN8 N$10 ADD_ONE GND GND n L=2u W=6u
        MP505 N$12429 N$12633 VDD VDD p L=2u W=6u
        MN505 N$12429 N$12633 GND GND n L=2u W=6u
        MN404 N$1177 GND GND GND n L=2u W=5u
        MN591 SK3 N$1491 GND GND n L=2u W=6u
        MP502 N$1571 N$1570 VDD VDD p L=2u W=6u
        MP517 N$1559 N$1558 VDD VDD p L=2u W=5u
        MP518 N$1557 N$11083 N$1559 VDD p L=2u W=5u
        MN267 N$310 N$311 GND GND n L=2u W=6u
        MP267 N$310 N$311 VDD VDD p L=2u W=6u
        MP61 N$271 CK N$282 VDD p L=2u W=6u
        MP269 N$306 CK VDD VDD p L=2u W=5u
        MN748 N$11332 N$11333 N$11083 GND n L=2u W=6u
        MN403 N$1177 N$1179 GND GND n L=2u W=5u
        MN268 N$311 N$309 GND GND n L=2u W=6u
        MP268 N$311 N$309 VDD VDD p L=2u W=6u
        MP450 N$1619 N$1620 N$1622 VDD p L=2u W=3u
        MP8 N$10 ADD_ONE VDD VDD p L=2u W=6u
        MN369 N$394 N$409 N$397 GND n L=2u W=5u
        MP333 N$345 N$11347 N$14091 VDD p L=2u W=5u
        MN326 N$14091 N$11347 GND GND n L=2u W=5u
        MP370 GND N$409 N$395 VDD p L=2u W=5u
        MN348 N$412 N$11347 N$331 GND n L=2u W=5u
        MP334 OUT8 N$11347 N$398 VDD p L=2u W=5u
        MP311 N$344 CK N$345 VDD p L=2u W=6u
        MN311 N$345 N$341 N$344 GND n L=2u W=6u
        MP310 N$342 N$341 N$344 VDD p L=2u W=6u
        MP252 N$242 CK N$298 VDD p L=2u W=6u
        MP254 N$301 N$298 VDD VDD p L=2u W=6u
        MP196 N$222 N$207 N$219 VDD p L=2u W=3u
        MN252 N$298 N$299 N$242 GND n L=2u W=6u
        MN150 N$166 N$162 GND GND n L=2u W=3u
        MP150 N$166 N$162 VDD VDD p L=2u W=3u
        MN149 N$162 N$138 N$164 GND n L=2u W=3u
        MN148 N$162 N$154 N$163 GND n L=2u W=3u
        MN117 N$127 N$102 GND GND n L=2u W=3u
        MN116 N$127 N$387 GND GND n L=2u W=3u
        MN308 N$343 N$340 GND GND n L=2u W=6u
        MP106 N$108 N$84 N$107 VDD p L=2u W=3u
        MP105 N$107 N$386 N$106 VDD p L=2u W=3u
        MP104 N$106 GND N$105 VDD p L=2u W=3u
        MP103 N$105 N$386 VDD VDD p L=2u W=3u
        MP102 N$105 GND VDD VDD p L=2u W=3u
        MP146 N$160 GND N$159 VDD p L=2u W=3u
        MP145 N$159 N$389 VDD VDD p L=2u W=3u
        MP144 N$159 GND VDD VDD p L=2u W=3u
        MP143 N$159 N$138 VDD VDD p L=2u W=3u
        MP187 N$210 N$394 VDD VDD p L=2u W=3u
        MP253 N$298 N$299 N$300 VDD p L=2u W=6u
        MN253 N$300 CK N$298 GND n L=2u W=6u
        MP294 N$331 N$332 VDD VDD p L=2u W=6u
        MP293 N$330 CK N$331 VDD p L=2u W=6u
        MN293 N$331 N$327 N$330 GND n L=2u W=6u
        MP292 N$328 N$327 N$330 VDD p L=2u W=6u
        MN292 N$330 CK N$328 GND n L=2u W=6u
        MN291 N$328 N$329 GND GND n L=2u W=6u
        MP345 N$14088 N$11347 N$376 VDD p L=2u W=5u
        MN344 N$411 N$11347 N$317 GND n L=2u W=5u
        MN13 N$20 N$21 N$23 GND n L=2u W=6u
        MP16 N$20 N$17 N$19 VDD p L=2u W=6u
        MP356 P1 N$409 N$386 VDD p L=2u W=5u
        MN402 N$11805 N$11794 GND GND n L=2u W=3u
        MN391 N$11570 N$13243 IN7 GND n L=2u W=5u
        MP391 IN7 N$13447 N$11570 VDD p L=2u W=5u
        MN390 N$11570 N$13447 N$1674 GND n L=2u W=5u
        MP390 N$1674 N$13243 N$11570 VDD p L=2u W=5u
        MN768 N$11802 N$11796 N$11803 GND n L=2u W=3u
        MN773 N$1599 N$11813 N$12429 GND n L=2u W=5u
        MN294 N$331 N$332 GND GND n L=2u W=6u
        MP773 N$12429 RST N$1599 VDD p L=2u W=5u
        MN772 N$1599 RST GND GND n L=2u W=5u
        MP772 GND N$11813 N$1599 VDD p L=2u W=5u
        MN771 N$11794 B0 GND GND n L=2u W=3u
        MP771 N$11794 B0 VDD VDD p L=2u W=3u
        MN485 N$1583 CK N$1585 GND n L=2u W=6u
        MN484 N$1585 N$1584 GND GND n L=2u W=6u
        MN354 N$385 N$409 N$398 GND n L=2u W=5u
        MP354 N$398 N$14096 N$385 VDD p L=2u W=5u
        MN353 N$385 N$14096 GND GND n L=2u W=5u
        MN343 N$411 N$14095 N$14087 GND n L=2u W=5u
        MP165 N$185 N$14079 VDD VDD p L=2u W=3u
        MP166 N$185 N$392 VDD VDD p L=2u W=3u
        MN313 N$346 N$344 GND GND n L=2u W=6u
        MP314 N$341 CK VDD VDD p L=2u W=5u
        MP98 N$100 N$84 N$96 VDD p L=2u W=3u
        MN345 N$376 N$14095 N$14088 GND n L=2u W=5u
        MN371 N$395 N$409 N$396 GND n L=2u W=5u
        MN305 N$334 CK GND GND n L=2u W=5u
        MP305 N$334 CK VDD VDD p L=2u W=5u
        MN304 N$339 N$337 GND GND n L=2u W=6u
        MN314 N$341 CK GND GND n L=2u W=5u
        MN98 N$104 N$386 GND GND n L=2u W=3u
        MN127 N$139 N$388 GND GND n L=2u W=3u
        MN126 N$140 N$388 GND GND n L=2u W=3u
        MN125 N$136 N$120 N$139 GND n L=2u W=3u
        MN124 N$139 GND GND GND n L=2u W=3u
        MN153 N$171 N$156 N$174 GND n L=2u W=3u
        MN152 N$174 N$14078 GND GND n L=2u W=3u
        MN151 N$173 N$171 GND GND n L=2u W=3u
        MP155 N$171 N$14078 N$170 VDD p L=2u W=3u
        MP154 N$171 N$156 N$168 VDD p L=2u W=3u
        MP123 N$132 GND VDD VDD p L=2u W=3u
        MP285 N$324 N$325 VDD VDD p L=2u W=6u
        MP284 N$323 CK N$324 VDD p L=2u W=6u
        MN284 N$324 N$320 N$323 GND n L=2u W=6u
        MP62 N$282 N$283 N$286 VDD p L=2u W=6u
        MN62 N$286 CK N$282 GND n L=2u W=6u
        MN66 N$361 N$283 N$288 GND n L=2u W=6u
        MP180 N$202 N$394 VDD VDD p L=2u W=3u
        MP179 N$202 N$14080 VDD VDD p L=2u W=3u
        MN285 N$324 N$325 GND GND n L=2u W=6u
        MN178 N$200 N$196 GND GND n L=2u W=3u
        MP178 N$200 N$196 VDD VDD p L=2u W=3u
        MN132 N$146 GND N$147 GND n L=2u W=3u
        MN131 N$145 N$120 GND GND n L=2u W=3u
        MP107 N$108 N$100 N$105 VDD p L=2u W=3u
        MN129 N$145 GND GND GND n L=2u W=3u
        MP135 N$144 N$136 N$141 VDD p L=2u W=3u
        MP134 N$144 N$120 N$143 VDD p L=2u W=3u
        MP133 N$143 N$388 N$142 VDD p L=2u W=3u
        MP132 N$142 GND N$141 VDD p L=2u W=3u
        MP176 N$196 N$173 N$195 VDD p L=2u W=3u
        MP175 N$195 N$392 N$194 VDD p L=2u W=3u
        MP174 N$194 N$14079 N$193 VDD p L=2u W=3u
        MP173 N$193 N$392 VDD VDD p L=2u W=3u
        MP202 N$228 N$14081 N$227 VDD p L=2u W=3u
        MP65 N$286 N$283 N$288 VDD p L=2u W=6u
        MP286 N$325 N$323 VDD VDD p L=2u W=6u
        MN254 N$301 N$298 GND GND n L=2u W=6u
        MN302 N$338 N$334 N$337 GND n L=2u W=6u
        MP301 N$335 N$334 N$337 VDD p L=2u W=6u
        MN301 N$337 CK N$335 GND n L=2u W=6u
        MN300 N$335 N$336 GND GND n L=2u W=6u
        MP300 N$335 N$336 VDD VDD p L=2u W=6u
        MN251 N$292 CK GND GND n L=2u W=5u
        MP251 N$292 CK VDD VDD p L=2u W=5u
        MN232 N$271 N$265 N$112 GND n L=2u W=5u
        MP195 N$221 N$395 N$219 VDD p L=2u W=3u
        MP194 N$219 N$395 VDD VDD p L=2u W=3u
        MP193 N$219 N$14081 VDD VDD p L=2u W=3u
        MP255 N$300 N$301 VDD VDD p L=2u W=6u
        MN192 N$217 N$213 GND GND n L=2u W=3u
        MN147 N$165 N$389 GND GND n L=2u W=3u
        MN146 N$164 GND N$165 GND n L=2u W=3u
        MN115 N$127 GND GND GND n L=2u W=3u
        MN144 N$163 N$389 GND GND n L=2u W=3u
        MN143 N$163 GND GND GND n L=2u W=3u
        MP149 N$162 N$154 N$159 VDD p L=2u W=3u
        MP148 N$162 N$138 N$161 VDD p L=2u W=3u
        MP147 N$161 N$389 N$160 VDD p L=2u W=3u
        MN199 N$231 N$14081 GND GND n L=2u W=3u
        MP205 N$230 N$222 N$227 VDD p L=2u W=3u
        MP204 N$230 N$207 N$229 VDD p L=2u W=3u
        MP203 N$229 N$395 N$228 VDD p L=2u W=3u
        MP225 N$217 N$265 N$262 VDD p L=2u W=5u
        MP67 N$361 N$290 VDD VDD p L=2u W=6u
        MP66 N$288 CK N$361 VDD p L=2u W=6u
        MP207 N$112 N$265 N$237 VDD p L=2u W=5u
        MN710 N$1385 N$1388 GND GND n L=2u W=6u
        MN177 N$196 N$173 N$198 GND n L=2u W=3u
        MP713 N$1384 CK N$14092 VDD p L=2u W=6u
        MN716 N$1387 CK GND GND n L=2u W=5u
        MP686 N$1402 CK N$14046 VDD p L=2u W=6u
        MN686 N$14046 N$14098 N$1402 GND n L=2u W=6u
        MP685 N$1404 N$14098 N$1402 VDD p L=2u W=6u
        MN685 N$1402 CK N$1404 GND n L=2u W=6u
        MN691 N$1398 CK N$1400 GND n L=2u W=6u
        MP690 N$1410 CK N$1400 VDD p L=2u W=6u
        MN690 N$1400 N$1399 N$1410 GND n L=2u W=6u
        MN689 N$14098 CK GND GND n L=2u W=5u
        MP689 N$14098 CK VDD VDD p L=2u W=5u
        MP644 N$1437 N$1441 VDD VDD p L=2u W=3u
        MN643 N$1441 N$1462 N$1439 GND n L=2u W=3u
        MN642 N$1441 N$1448 N$1440 GND n L=2u W=3u
        MN641 N$1438 N$1450 GND GND n L=2u W=3u
        MN647 N$1433 N$1447 N$1431 GND n L=2u W=3u
        MN646 N$1431 B3 GND GND n L=2u W=3u
        MN675 N$1410 N$1557 N$1452 GND n L=2u W=5u
        MP681 N$14097 CK N$1406 VDD p L=2u W=6u
        MN681 N$1406 N$14098 N$14097 GND n L=2u W=6u
        MN680 N$1408 N$1413 GND GND n L=2u W=5u
        MP680 GND N$1557 N$1408 VDD p L=2u W=5u
        MN679 N$1408 N$1557 N$1422 GND n L=2u W=5u
        MN880 N$14035 N$14040 GND GND n L=2u W=5u
        MP880 GND N$14037 N$14035 VDD p L=2u W=5u
        MN879 N$14035 N$14037 GND GND n L=2u W=5u
        MP879 GND N$14040 N$14035 VDD p L=2u W=5u
        MN878 N$14037 N$14040 GND GND n L=2u W=5u
        MP884 GND N$14037 N$14031 VDD p L=2u W=5u
        MN883 N$14031 N$14037 GND GND n L=2u W=5u
        MP883 GND N$14040 N$14031 VDD p L=2u W=5u
        MN882 N$14033 N$14040 GND GND n L=2u W=5u
        MP850 N$13966 N$14005 N$13965 VDD p L=2u W=3u
        MP849 N$13965 N$14005 VDD VDD p L=2u W=3u
        MP848 N$13965 N$14090 VDD VDD p L=2u W=3u
        MN847 OUT5 N$13959 GND GND n L=2u W=3u
        MN875 OUT7 N$13991 GND GND n L=2u W=3u
        MP875 OUT7 N$13991 VDD VDD p L=2u W=3u
        MN874 N$13991 N$13969 N$13993 GND n L=2u W=3u
        MN873 N$13991 N$13983 N$13992 GND n L=2u W=3u
        MP160 N$177 N$14078 N$176 VDD p L=2u W=3u
        MP159 N$176 N$390 VDD VDD p L=2u W=3u
        MN751 N$11334 N$11335 GND GND n L=2u W=6u
        MP751 N$11334 N$11335 VDD VDD p L=2u W=6u
        MN750 N$11335 N$11332 GND GND n L=2u W=6u
        MN736 N$11328 CK N$11326 GND n L=2u W=6u
        MP735 N$11344 CK N$11326 VDD p L=2u W=6u
        MN735 N$11326 N$11327 N$11344 GND n L=2u W=6u
        MN734 N$11321 CK GND GND n L=2u W=5u
        MP734 N$11321 CK VDD VDD p L=2u W=5u
        MN733 N$11325 N$11324 GND GND n L=2u W=6u
        MP733 N$11325 N$11324 VDD VDD p L=2u W=6u
        MN732 N$11099 N$11325 GND GND n L=2u W=6u
        MP353 GND N$409 N$385 VDD p L=2u W=5u
        MP359 N$410 N$14096 N$387 VDD p L=2u W=5u
        MN359 N$387 N$409 N$410 GND n L=2u W=5u
        MP360 P3 N$409 N$388 VDD p L=2u W=5u
        MN360 N$388 N$14096 P3 GND n L=2u W=5u
        MN164 N$183 N$179 GND GND n L=2u W=3u
        MP164 N$183 N$179 VDD VDD p L=2u W=3u
        MN163 N$179 N$156 N$181 GND n L=2u W=3u
        MN162 N$179 N$171 N$180 GND n L=2u W=3u
        MN295 N$332 N$330 GND GND n L=2u W=6u
        MP161 N$178 N$390 N$177 VDD p L=2u W=3u
        MP113 N$118 GND N$117 VDD p L=2u W=3u
        MP112 N$118 N$102 N$114 VDD p L=2u W=3u
        MP111 N$117 N$387 N$114 VDD p L=2u W=3u



*.ends mynand3

* Auxiliary circuit for power analysis
Cp Pav 0 100p
Rp Pav 0 100k
Fp 0 Pav Vtstp 0.003125
*Output load capacitance if you have any

*Cload1 out GND 200fF
.MODEL n NMOS LEVEL = 3
+ TOX = 200E-10 NSUB = 1E17 GAMMA = 0.5
+ PHI = 0.7 VTO = 0.8 DELTA = 3.0
+ UO = 650 ETA = 3.0E-6 THETA = 0.1
+ KP = 120E-6 VMAX = 1E5 KAPPA = 0.3
+ RSH = 0 NFS = 1E12 TPG = 1
+ XJ = 500E-9 LD = 100E-9
+ CGDO = 200E-12 CGSO = 200E-12 CGBO = 1E-10
+ CJ = 400E-6 PB = 1 MJ = 0.5
+ CJSW = 300E-12 MJSW = 0.5

.MODEL p PMOS LEVEL = 3
+ TOX = 200E-10 NSUB = 1E17 GAMMA = 0.6
+ PHI = 0.7 VTO = -0.9 DELTA = 0.1
+ UO = 250 ETA = 0 THETA = 0.1
+ KP = 40E-6 VMAX = 5E4 KAPPA = 1
+ RSH = 0 NFS = 1E12 TPG = -1
+ XJ = 500E-9 LD = 100E-9
+ CGDO = 200E-12 CGSO = 200E-12 CGBO = 1E-10
+ CJ = 400E-6 PB = 1 MJ = 0.5
+ CJSW = 300E-12 MJSW = 0.5

*Define power rails
Vddt top 0 5
Vtstp top Vdd 0
Vss GND 0 0

* Define input voltages of A and B

Vck CK 0 PWL(0 5 20N 5 20.1N 0 40N 0 40.1N 5 60N 5 60.1N 0 80N 0 80.1N 5 100N 5 
+ 100.1N 0 120N 0 120.1N 5 140N 5 140.1N 0 160N 0 160.1N 5 180N 5 180.1N 0 200N 0
+ 200.1N 5 220N 5 220.1N 0 240N 0 240.1N 5 260N 5 260.1N 0 280N 0 280.1N 5 300N 5 
+ 300.1N 0 320N 0 320.1N 5 340N 5 340.1N 0 360N 0 360.1N 5 380N 5 380.1N 0 400N 0 
+ 400.1N 5 420N 5 420.1N 0 440N 0 440.1N 5 460N 5 460.1N 0 480N 0 480.1N 5 500N 5)

Va5 A5 0 PWL(0 5 20N 5 20.1N 5 40N 5 40.1N 5 60N 5 60.1N 5 80N 5 80.1N 5 100N 5 
+ 100.1N 5 120N 5 120.1N 5 140N 5 140.1N 5 160N 5 160.1N 5 180N 5 180.1N 5 200N 5
+ 200.1N 0 220N 0 220.1N 0 240N 0 240.1N 0 260N 0 260.1N 0 280N 0 280.1N 0 300N 0 
+ 300.1N 0 320N 0 320.1N 0 340N 0 340.1N 0 360N 0 360.1N 0 380N 0 380.1N 0 400N 0 
+ 400.1N 0 420N 0 420.1N 0 440N 0 440.1N 0 460N 0 460.1N 0 480N 0 480.1N 0 500N 0)

Vp1 P1 0 PWL(0 5 20N 5 20.1N 5 40N 5 40.1N 5 60N 5 60.1N 5 80N 5 80.1N 5 100N 5 
+ 100.1N 5 120N 5 120.1N 5 140N 5 140.1N 5 160N 5 160.1N 5 180N 5 180.1N 5 200N 5
+ 200.1N 5 220N 5 220.1N 5 240N 5 240.1N 5 260N 5 260.1N 5 280N 5 280.1N 5 300N 5 
+ 300.1N 5 320N 5 320.1N 5 340N 5 340.1N 5 360N 5 360.1N 5 380N 5 380.1N 5 400N 5 
+ 400.1N 5 420N 5 420.1N 5 440N 5 440.1N 5 460N 5 460.1N 5 480N 5 480.1N 5 500N 5)


Vp2 P2 0 PWL(0 0 20N 0 20.1N 0 40N 0 40.1N 0 60N 0 60.1N 0 80N 0 80.1N 0 100N 0 
+ 100.1N 0 120N 0 120.1N 0 140N 0 140.1N 0 160N 0 160.1N 0 180N 0 180.1N 0 200N 0
+ 200.1N 0 220N 0 220.1N 0 240N 0 240.1N 0 260N 0 260.1N 0 280N 0 280.1N 0 300N 0 
+ 300.1N 0 320N 0 320.1N 0 340N 0 340.1N 0 360N 0 360.1N 0 380N 0 380.1N 0 400N 0 
+ 400.1N 0 420N 0 420.1N 0 440N 0 440.1N 0 460N 0 460.1N 0 480N 0 480.1N 0 500N 0)

Vp3 P3 0 PWL(0 5 20N 5 20.1N 5 40N 5 40.1N 5 60N 5 60.1N 5 80N 5 80.1N 5 100N 5 
+ 100.1N 5 120N 5 120.1N 5 140N 5 140.1N 5 160N 5 160.1N 5 180N 5 180.1N 5 200N 5
+ 200.1N 5 220N 5 220.1N 5 240N 5 240.1N 5 260N 5 260.1N 5 280N 5 280.1N 5 300N 5 
+ 300.1N 5 320N 5 320.1N 5 340N 5 340.1N 5 360N 5 360.1N 5 380N 5 380.1N 5 400N 5 
+ 400.1N 5 420N 5 420.1N 5 440N 5 440.1N 5 460N 5 460.1N 5 480N 5 480.1N 5 500N 5)


Vp4 P4 0 PWL(0 0 20N 0 20.1N 0 40N 0 40.1N 0 60N 0 60.1N 0 80N 0 80.1N 0 100N 0 
+ 100.1N 0 120N 0 120.1N 0 140N 0 140.1N 0 160N 0 160.1N 0 180N 0 180.1N 0 200N 0
+ 200.1N 0 220N 0 220.1N 0 240N 0 240.1N 0 260N 0 260.1N 0 280N 0 280.1N 0 300N 0 
+ 300.1N 0 320N 0 320.1N 0 340N 0 340.1N 0 360N 0 360.1N 0 380N 0 380.1N 0 400N 0 
+ 400.1N 0 420N 0 420.1N 0 440N 0 440.1N 0 460N 0 460.1N 0 480N 0 480.1N 0 500N 0)

Vrst RST 0 PWL(0 5 20N 5 20.1N 5 40N 5 40.1N 0 60N 0 60.1N 0 80N 0 80.1N 0 100N 0 
+ 100.1N 0 120N 0 120.1N 0 140N 0 140.1N 0 160N 0 160.1N 0 180N 0 180.1N 0 200N 0
+ 200.1N 0 220N 0 220.1N 0 240N 0 240.1N 0 260N 0 260.1N 0 280N 0 280.1N 0 300N 0 
+ 300.1N 0 320N 0 320.1N 0 340N 0 340.1N 0 360N 0 360.1N 0 380N 0 380.1N 0 400N 0 
+ 400.1N 0 420N 0 420.1N 0 440N 0 440.1N 0 460N 0 460.1N 0 480N 0 480.1N 0 500N 0)

Vb0 B0 0 PWL(0 5 20N 5 20.1N 5 40N 5 40.1N 5 60N 5 60.1N 5 80N 5 80.1N 5 100N 5 
+ 100.1N 5 120N 5 120.1N 5 140N 5 140.1N 5 160N 5 160.1N 5 180N 5 180.1N 5 200N 5
+ 200.1N 5 220N 5 220.1N 5 240N 5 240.1N 5 260N 5 260.1N 5 280N 5 280.1N 5 300N 5 
+ 300.1N 5 320N 5 320.1N 5 340N 5 340.1N 5 360N 5 360.1N 5 380N 5 380.1N 5 400N 5 
+ 400.1N 5 420N 5 420.1N 5 440N 5 440.1N 5 460N 5 460.1N 5 480N 5 480.1N 5 500N 5)

Vb1 B1 0 PWL(0 0 20N 0 20.1N 0 40N 0 40.1N 0 60N 0 60.1N 0 80N 0 80.1N 0 100N 0 
+ 100.1N 0 120N 0 120.1N 0 140N 0 140.1N 0 160N 0 160.1N 0 180N 0 180.1N 0 200N 0
+ 200.1N 0 220N 0 220.1N 0 240N 0 240.1N 0 260N 0 260.1N 0 280N 0 280.1N 0 300N 0 
+ 300.1N 0 320N 0 320.1N 0 340N 0 340.1N 0 360N 0 360.1N 0 380N 0 380.1N 0 400N 0 
+ 400.1N 0 420N 0 420.1N 0 440N 0 440.1N 0 460N 0 460.1N 0 480N 0 480.1N 0 500N 0)

Vb2 B2 0 PWL(0 5 20N 5 20.1N 5 40N 5 40.1N 5 60N 5 60.1N 5 80N 5 80.1N 5 100N 5 
+ 100.1N 5 120N 5 120.1N 5 140N 5 140.1N 5 160N 5 160.1N 5 180N 5 180.1N 5 200N 5
+ 200.1N 5 220N 5 220.1N 5 240N 5 240.1N 5 260N 5 260.1N 5 280N 5 280.1N 5 300N 5 
+ 300.1N 5 320N 5 320.1N 5 340N 5 340.1N 5 360N 5 360.1N 5 380N 5 380.1N 5 400N 5 
+ 400.1N 5 420N 5 420.1N 5 440N 5 440.1N 5 460N 5 460.1N 5 480N 5 480.1N 5 500N 5)

Vb3 B3 0 PWL(0 0 20N 0 20.1N 0 40N 0 40.1N 0 60N 0 60.1N 0 80N 0 80.1N 0 100N 0 
+ 100.1N 0 120N 0 120.1N 0 140N 0 140.1N 0 160N 0 160.1N 0 180N 0 180.1N 0 200N 0
+ 200.1N 0 220N 0 220.1N 0 240N 0 240.1N 0 260N 0 260.1N 0 280N 0 280.1N 0 300N 0 
+ 300.1N 0 320N 0 320.1N 0 340N 0 340.1N 0 360N 0 360.1N 0 380N 0 380.1N 0 400N 0 
+ 400.1N 0 420N 0 420.1N 0 440N 0 440.1N 0 460N 0 460.1N 0 480N 0 480.1N 0 500N 0)

Vc C 0 PWL(0 5 20N 5 20.1N 5 40N 5 40.1N 5 60N 5 60.1N 5 80N 5 80.1N 5 100N 5 
+ 100.1N 5 120N 5 120.1N 5 140N 5 140.1N 5 160N 5 160.1N 5 180N 5 180.1N 5 200N 5
+ 200.1N 5 220N 5 220.1N 5 240N 5 240.1N 5 260N 5 260.1N 5 280N 5 280.1N 5 300N 5 
+ 300.1N 5 320N 5 320.1N 5 340N 5 340.1N 5 360N 5 360.1N 5 380N 5 380.1N 5 400N 5 
+ 400.1N 5 420N 5 420.1N 5 440N 5 440.1N 5 460N 5 460.1N 5 480N 5 480.1N 5 500N 5)

Vadd_one add_one 0 PWL(0 5 20N 5 20.1N 5 40N 5 40.1N 5 60N 5 60.1N 5 80N 5 80.1N 5 100N 5 
+ 100.1N 5 120N 5 120.1N 5 140N 5 140.1N 5 160N 5 160.1N 5 180N 5 180.1N 5 200N 5
+ 200.1N 5 220N 5 220.1N 5 240N 5 240.1N 5 260N 5 260.1N 5 280N 5 280.1N 5 300N 5 
+ 300.1N 5 320N 5 320.1N 5 340N 5 340.1N 5 360N 5 360.1N 5 380N 5 380.1N 5 400N 5 
+ 400.1N 5 420N 5 420.1N 5 440N 5 440.1N 5 460N 5 460.1N 5 480N 5 480.1N 5 500N 5)


*Define transient simulation and probe voltage/current signals
.TRAN 20N 500N
.PROBE V(*) I(*)
.end
