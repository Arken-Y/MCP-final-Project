




*.subckt mynand3 A B GND Out Vdd



* MAIN CELL: Component pathname : /home/mentor/jack/jaggu
*
               MP605 N$8587 N$8586 N$8585 VDD p L=2u W=3u
        MN642 N$6397 N$6404 N$6396 GND n L=2u W=3u
        MP636 N$6403 N$6404 VDD VDD p L=2u W=3u
        MP637 N$6400 N$6418 VDD VDD p L=2u W=3u
        MP642 N$6397 N$6418 N$6398 VDD p L=2u W=3u
        MP640 N$6399 H2 N$6400 VDD p L=2u W=3u
        MP641 N$6398 N$6406 N$6399 VDD p L=2u W=3u
        MP621 N$6419 H1 N$6420 VDD p L=2u W=3u
        MP620 N$6419 N$8383 N$6422 VDD p L=2u W=3u
        MP619 N$6420 N$6421 N$6422 VDD p L=2u W=3u
        MP618 N$6422 N$6421 VDD VDD p L=2u W=3u
        MP617 N$6422 H1 VDD VDD p L=2u W=3u
        MN635 N$6402 N$6406 GND GND n L=2u W=3u
        MN636 N$6404 H2 N$6401 GND n L=2u W=3u
        MN622 N$6419 H1 N$6416 GND n L=2u W=3u
        MN621 N$6417 N$6421 GND GND n L=2u W=3u
        MP604 N$8585 N$8586 VDD VDD p L=2u W=3u
        MP603 N$8585 H0 VDD VDD p L=2u W=3u
        MP679 N$6378 N$6376 N$6368 VDD p L=2u W=5u
        MN684 N$6364 N$6363 GND GND n L=2u W=6u
        MP651 N$6385 N$6403 VDD VDD p L=2u W=3u
        MN656 N$6382 N$6389 N$6381 GND n L=2u W=3u
        MN655 N$6379 N$6391 GND GND n L=2u W=3u
        MN654 N$6380 H3 N$6379 GND n L=2u W=3u
        MN682 N$6364 CK N$6366 GND n L=2u W=6u
        MN687 N$6268 N$6361 GND GND n L=2u W=6u
        MP687 N$6268 N$6361 VDD VDD p L=2u W=6u
        MP660 N$6421 N$6444 VDD VDD p L=2u W=3u
        MN679 N$6368 N$6515 N$6378 GND n L=2u W=5u
        MP680 GND N$6515 N$6368 VDD p L=2u W=5u
        MN685 N$6362 CK N$6364 GND n L=2u W=6u
        MN551 N$6488 N$6499 GND GND n L=2u W=5u
        MP551 N$6488 N$6499 VDD VDD p L=2u W=5u
        MN556 N$6483 N$6499 N$6490 GND n L=2u W=5u
        MP556 N$6490 N$6488 N$6483 VDD p L=2u W=5u
        MN555 N$6484 N$6488 GND GND n L=2u W=5u
        MP555 GND N$6499 N$6484 VDD p L=2u W=5u
        MN554 N$6484 N$6499 N$6526 GND n L=2u W=5u
        MP554 N$6526 N$6488 N$6484 VDD p L=2u W=5u
        MP559 N$6481 N$6480 N$6477 VDD p L=2u W=6u
        MN559 N$6477 CK N$6481 GND n L=2u W=6u
        MP558 N$6479 CK N$6481 VDD p L=2u W=6u
        MN558 N$6481 N$6480 N$6479 GND n L=2u W=6u
        MN557 N$6483 N$6488 GND GND n L=2u W=5u
        MP557 GND N$6499 N$6483 VDD p L=2u W=5u
        MN609 N$8595 H0 GND GND n L=2u W=3u
        MP207 GND N$7766 N$6919 VDD p L=2u W=5u
        MN206 N$6920 N$7766 GND GND n L=2u W=5u
        MP206 GND N$6904 N$6920 VDD p L=2u W=5u
        MN569 N$6468 N$6472 GND GND n L=2u W=6u
        MP575 N$6471 CK VDD VDD p L=2u W=5u
        MN574 N$6465 N$6467 GND GND n L=2u W=6u
        MP217 N$6714 N$6910 N$6730 VDD p L=2u W=5u
        MP225 N$6918 N$6905 N$6914 VDD p L=2u W=5u
        MP572 N$6467 CK N$6910 VDD p L=2u W=6u
        MP578 N$6460 N$6464 VDD VDD p L=2u W=6u
        MP577 N$6464 N$6463 N$6461 VDD p L=2u W=6u
        MN577 N$6461 CK N$6464 GND n L=2u W=6u
        MP576 N$6462 CK N$6464 VDD p L=2u W=6u
        MP241 N$6944 N$6911 N$6895 VDD p L=2u W=5u
        MP351 N$6948 N$6913 N$6895 VDD p L=2u W=5u
        MN240 N$6894 N$6911 N$6914 GND n L=2u W=5u
        MP240 N$6914 N$6913 N$6894 VDD p L=2u W=5u
        MN239 N$6894 N$6913 N$6732 GND n L=2u W=5u
        MP239 N$6732 N$6911 N$6894 VDD p L=2u W=5u
        MN241 N$6895 N$6913 N$6944 GND n L=2u W=5u
        MN238 N$6913 N$6911 GND GND n L=2u W=5u
        MP238 N$6913 N$6911 VDD VDD p L=2u W=5u
        MP352 N$6914 N$6911 N$6896 VDD p L=2u W=5u
        MN237 N$6893 N$6911 N$6944 GND n L=2u W=5u
        MP237 N$6944 N$6913 N$6893 VDD p L=2u W=5u
        MN234 N$6893 N$6913 N$6730 GND n L=2u W=5u
        MP234 N$6730 N$6911 N$6893 VDD p L=2u W=5u
        MN233 N$6945 N$6910 GND GND n L=2u W=5u
        MP233 GND N$6905 N$6945 VDD p L=2u W=5u
        MN659 N$8586 N$9213 GND GND n L=2u W=3u
        MP659 N$8586 N$9213 VDD VDD p L=2u W=3u
        MN616 N$9216 N$8594 GND GND n L=2u W=3u
        MN617 N$6418 N$6419 GND GND n L=2u W=3u
        MN560 N$6476 N$6481 GND GND n L=2u W=6u
        MP560 N$6476 N$6481 VDD VDD p L=2u W=6u
        MP566 N$6480 CK VDD VDD p L=2u W=5u
        MN565 N$6473 N$6475 GND GND n L=2u W=6u
        MP624 N$6415 H1 VDD VDD p L=2u W=3u
        MP623 N$6415 N$8383 VDD VDD p L=2u W=3u
        MP622 N$6418 N$6419 VDD VDD p L=2u W=3u
        MP563 N$6475 CK HK_SK VDD p L=2u W=6u
        MN563 HK_SK N$6480 N$6475 GND n L=2u W=6u
        MP569 N$6468 N$6472 VDD VDD p L=2u W=6u
        MN624 N$6411 N$6421 GND GND n L=2u W=3u
        MP594 N$6533 N$6447 N$9213 VDD p L=2u W=5u
        MN226 N$6948 N$6905 N$6918 GND n L=2u W=5u
        MP226 N$6918 N$6910 N$6948 VDD p L=2u W=5u
        MN378 N$6955 N$6911 GND GND n L=2u W=5u
        MP378 GND N$6913 N$6955 VDD p L=2u W=5u
        MN377 N$6955 N$6913 N$6945 GND n L=2u W=5u
        MP377 N$6945 N$6911 N$6955 VDD p L=2u W=5u
        MP383 N$6747 N$6221 N$6746 VDD p L=2u W=3u
        MN376 N$6956 N$6911 GND GND n L=2u W=5u
        MP376 GND N$6913 N$6956 VDD p L=2u W=5u
        MN375 N$6956 N$6913 N$6946 GND n L=2u W=5u
        MP375 N$6946 N$6911 N$6956 VDD p L=2u W=5u
        MP382 N$6747 GND N$6745 VDD p L=2u W=3u
        MN374 N$6957 N$6911 N$6945 GND n L=2u W=5u
        MP374 N$6945 N$6913 N$6957 VDD p L=2u W=5u
        MN373 N$6957 N$6913 N$6947 GND n L=2u W=5u
        MP373 N$6947 N$6911 N$6957 VDD p L=2u W=5u
        MN371 N$6883 N$6913 N$6948 GND n L=2u W=5u
        MN372 N$6883 N$6911 N$6946 GND n L=2u W=5u
        MP372 N$6946 N$6913 N$6883 VDD p L=2u W=5u
        MP381 N$6746 N$6900 N$6745 VDD p L=2u W=3u
        MP585 N$6454 CK N$6456 VDD p L=2u W=6u
        MN585 N$6456 N$6455 N$6454 GND n L=2u W=6u
        MP590 N$6451 CK S3 VDD p L=2u W=6u
        MN590 S3 N$6455 N$6451 GND n L=2u W=6u
        MP230 N$6916 N$6910 N$6946 VDD p L=2u W=5u
        MN229 N$6947 N$6910 N$6916 GND n L=2u W=5u
        MP229 N$6916 N$6905 N$6947 VDD p L=2u W=5u
        MN225 N$6914 N$6910 N$6918 GND n L=2u W=5u
        MN216 N$6915 N$7766 GND GND n L=2u W=5u
        MP216 GND N$6904 N$6915 VDD p L=2u W=5u
        MN215 N$6915 N$6904 A0 GND n L=2u W=5u
        MN584 N$6463 CK GND GND n L=2u W=5u
        MP593 N$6455 CK VDD VDD p L=2u W=5u
        MN592 N$6449 N$6451 GND GND n L=2u W=6u
        MP592 N$6449 N$6451 VDD VDD p L=2u W=6u
        MN591 S3 N$6449 GND GND n L=2u W=6u
        MP591 S3 N$6449 VDD VDD p L=2u W=6u
        MN596 N$6447 N$6515 GND GND n L=2u W=5u
        MP596 N$6447 N$6515 VDD VDD p L=2u W=5u
        MN595 N$9213 N$6447 GND GND n L=2u W=5u
        MP595 GND N$6515 N$9213 VDD p L=2u W=5u
        MP224 N$6919 N$6910 N$6914 VDD p L=2u W=5u
        MN223 N$6944 N$6910 N$6919 GND n L=2u W=5u
        MP223 N$6919 N$6905 N$6944 VDD p L=2u W=5u
        MN222 N$6944 N$6905 N$6920 GND n L=2u W=5u
        MP222 N$6920 N$6910 N$6944 VDD p L=2u W=5u
        MN221 N$6732 N$6910 N$6920 GND n L=2u W=5u
        MP221 N$6920 N$6905 N$6732 VDD p L=2u W=5u
        MN220 N$6732 N$6905 N$6864 GND n L=2u W=5u
        MP220 N$6864 N$6910 N$6732 VDD p L=2u W=5u
        MN230 N$6946 N$6905 N$6916 GND n L=2u W=5u
        MP865 GND N$6884 N$6900 VDD p L=2u W=5u
        MN864 N$6900 N$6884 N$6955 GND n L=2u W=5u
        MP864 N$6955 S3 N$6900 VDD p L=2u W=5u
        MN863 N$6696 S3 GND GND n L=2u W=5u
        MP863 GND N$6884 N$6696 VDD p L=2u W=5u
        MN862 N$6696 N$6884 N$6956 GND n L=2u W=5u
        MP862 N$6956 S3 N$6696 VDD p L=2u W=5u
        MN861 N$6887 S3 GND GND n L=2u W=5u
        MP861 GND N$6884 N$6887 VDD p L=2u W=5u
        MN860 N$6887 N$6884 N$6957 GND n L=2u W=5u
        MN116 GND N$6688 N$6660 GND n L=2u W=5u
        MN115 N$6660 N$6328 A1 GND n L=2u W=5u
        MP116 N$6660 N$6328 GND VDD p L=2u W=5u
        MP115 A1 N$6688 N$6660 VDD p L=2u W=5u
        MN114 GND N$6687 N$6659 GND n L=2u W=5u
        MN113 N$6659 N$6685 A0 GND n L=2u W=5u
        MP114 N$6659 N$6685 GND VDD p L=2u W=5u
        MP113 A0 N$6687 N$6659 VDD p L=2u W=5u
        MP330 N$6169 N$8380 N$6931 VDD p L=2u W=5u
        MP120 N$6664 N$6691 GND VDD p L=2u W=5u
        MP119 A3 N$6319 N$6664 VDD p L=2u W=5u
        MN118 GND N$6692 N$6662 GND n L=2u W=5u
        MN117 N$6662 N$6690 A2 GND n L=2u W=5u
        MP118 N$6662 N$6690 GND VDD p L=2u W=5u
        MN232 N$6945 N$6905 N$6915 GND n L=2u W=5u
        MP232 N$6915 N$6910 N$6945 VDD p L=2u W=5u
        MN231 N$6946 N$6910 N$6915 GND n L=2u W=5u
        MP231 N$6915 N$6905 N$6946 VDD p L=2u W=5u
        MN336 N$6933 N$8380 GND GND n L=2u W=5u
        MP336 N$6933 N$8380 VDD VDD p L=2u W=5u
        MN335 N$6246 N$8380 N$6211 GND n L=2u W=5u
        MP204 GND N$6904 N$6864 VDD p L=2u W=5u
        MN203 N$6864 N$6904 GND GND n L=2u W=5u
        MP588 N$6453 N$6452 VDD VDD p L=2u W=6u
        MN593 N$6455 CK GND GND n L=2u W=5u
        MN797 N$6809 N$6889 GND GND n L=2u W=3u
        MN796 N$6810 N$6889 GND GND n L=2u W=3u
        MN795 N$6806 N$6793 N$6809 GND n L=2u W=3u
        MN794 N$6809 N$6924 GND GND n L=2u W=3u
        MN793 N$6808 N$6806 GND GND n L=2u W=3u
        MP797 N$6806 N$6924 N$6805 VDD p L=2u W=3u
        MP796 N$6806 N$6793 N$6804 VDD p L=2u W=3u
        MP795 N$6805 N$6889 N$6804 VDD p L=2u W=3u
        MP794 N$6804 N$6889 VDD VDD p L=2u W=3u
        MP793 N$6804 N$6924 VDD VDD p L=2u W=3u
        MN798 N$6806 N$6924 N$6810 GND n L=2u W=3u
        MN792 OUT3 N$6799 GND GND n L=2u W=3u
        MP792 OUT3 N$6799 VDD VDD p L=2u W=3u
        MN791 N$6799 N$6865 N$6801 GND n L=2u W=3u
        MN790 N$6799 N$6791 N$6800 GND n L=2u W=3u
        MN789 N$6802 N$6888 GND GND n L=2u W=3u
        MN788 N$6801 N$6923 N$6802 GND n L=2u W=3u
        MN787 N$6800 N$6865 GND GND n L=2u W=3u
        MN219 N$6905 N$6910 GND GND n L=2u W=5u
        MP219 N$6905 N$6910 VDD VDD p L=2u W=5u
        MN204 N$6864 N$7766 GND GND n L=2u W=5u
        MP789 N$6798 N$6888 N$6797 VDD p L=2u W=3u
        MP788 N$6797 N$6923 N$6796 VDD p L=2u W=3u
        MP787 N$6796 N$6888 VDD VDD p L=2u W=3u
        MP786 N$6796 N$6923 VDD VDD p L=2u W=3u
        MP850 N$6896 N$6884 N$6891 VDD p L=2u W=5u
        MN849 N$6891 N$6884 N$6893 GND n L=2u W=5u
        MP849 N$6893 S3 N$6891 VDD p L=2u W=5u
        MP831 N$6843 N$6890 N$6842 VDD p L=2u W=3u
        MP830 N$6842 N$6931 N$6841 VDD p L=2u W=3u
        MN848 OUT7 N$6858 GND GND n L=2u W=3u
        MP848 OUT7 N$6858 VDD VDD p L=2u W=3u
        MN847 N$6858 N$6838 N$6860 GND n L=2u W=3u
        MN846 N$6858 N$6851 N$6859 GND n L=2u W=3u
        MN845 N$6861 N$6891 GND GND n L=2u W=3u
        MN844 N$6860 N$6930 N$6861 GND n L=2u W=3u
        MN843 N$6859 N$6838 GND GND n L=2u W=3u
        MN842 N$6859 N$6891 GND GND n L=2u W=3u
        MN841 N$6859 N$6930 GND GND n L=2u W=3u
        MP847 N$6858 N$6851 N$6855 VDD p L=2u W=3u
        MP846 N$6858 N$6838 N$6857 VDD p L=2u W=3u
        MP567 N$6470 CK N$6472 VDD p L=2u W=6u
        MN567 N$6472 N$6471 N$6470 GND n L=2u W=6u
        MN566 N$6480 CK GND GND n L=2u W=5u
        MN594 N$9213 N$6515 N$6533 GND n L=2u W=5u
        MN572 N$6910 N$6471 N$6467 GND n L=2u W=6u
        MN786 N$6800 N$6888 GND GND n L=2u W=3u
        MN785 N$6800 N$6923 GND GND n L=2u W=3u
        MP791 N$6799 N$6791 N$6796 VDD p L=2u W=3u
        MP790 N$6799 N$6865 N$6798 VDD p L=2u W=3u
        MN310 N$6156 CK N$6158 GND n L=2u W=6u
        MN309 N$6158 N$6157 GND GND n L=2u W=6u
        MN314 N$6159 CK GND GND n L=2u W=5u
        MP785 N$6796 N$6865 VDD VDD p L=2u W=3u
        MP784 N$6793 N$6791 VDD VDD p L=2u W=3u
        MN784 N$6791 N$6923 N$6795 GND n L=2u W=3u
        MP815 N$6826 N$6867 VDD VDD p L=2u W=3u
        MP814 N$6826 N$6925 VDD VDD p L=2u W=3u
        MP845 N$6857 N$6891 N$6856 VDD p L=2u W=3u
        MP844 N$6856 N$6930 N$6855 VDD p L=2u W=3u
        MP843 N$6855 N$6891 VDD VDD p L=2u W=3u
        MP842 N$6855 N$6930 VDD VDD p L=2u W=3u
        MP841 N$6855 N$6838 VDD VDD p L=2u W=3u
        MP840 CARRY_OUT N$6851 VDD VDD p L=2u W=3u
        MN840 N$6851 N$6930 N$6854 GND n L=2u W=3u
        MN839 N$6853 N$6891 GND GND n L=2u W=3u
        MN838 N$6854 N$6891 GND GND n L=2u W=3u
        MN837 N$6851 N$6838 N$6853 GND n L=2u W=3u
        MN836 N$6853 N$6930 GND GND n L=2u W=3u
        MN835 CARRY_OUT N$6851 GND GND n L=2u W=3u
        MP839 N$6851 N$6930 N$6850 VDD p L=2u W=3u
        MP838 N$6851 N$6838 N$6849 VDD p L=2u W=3u
        MP837 N$6850 N$6891 N$6849 VDD p L=2u W=3u
        MP836 N$6849 N$6891 VDD VDD p L=2u W=3u
        MP835 N$6849 N$6930 VDD VDD p L=2u W=3u
        MN587 N$6452 N$6456 GND GND n L=2u W=6u
        MP587 N$6452 N$6456 VDD VDD p L=2u W=6u
        MP586 N$6456 N$6455 N$6453 VDD p L=2u W=6u
        MN586 N$6453 CK N$6456 GND n L=2u W=6u
        MN832 N$6844 N$6836 N$6845 GND n L=2u W=3u
        MN831 N$6847 N$6890 GND GND n L=2u W=3u
        MN830 N$6846 N$6931 N$6847 GND n L=2u W=3u
        MN829 N$6845 N$6823 GND GND n L=2u W=3u
        MP589 N$6453 N$6455 N$6451 VDD p L=2u W=6u
        MN589 N$6451 CK N$6453 GND n L=2u W=6u
        MN588 N$6453 N$6452 GND GND n L=2u W=6u
        MP832 N$6844 N$6823 N$6843 VDD p L=2u W=3u
        MP799 N$6811 N$6793 VDD VDD p L=2u W=3u
        MP798 N$6808 N$6806 VDD VDD p L=2u W=3u
        MP829 N$6841 N$6890 VDD VDD p L=2u W=3u
        MP828 N$6841 N$6931 VDD VDD p L=2u W=3u
        MP827 N$6841 N$6823 VDD VDD p L=2u W=3u
        MP826 N$6838 N$6836 VDD VDD p L=2u W=3u
        MN826 N$6836 N$6931 N$6840 GND n L=2u W=3u
        MN825 N$6839 N$6890 GND GND n L=2u W=3u
        MN824 N$6840 N$6890 GND GND n L=2u W=3u
        MN823 N$6836 N$6823 N$6839 GND n L=2u W=3u
        MN822 N$6839 N$6931 GND GND n L=2u W=3u
        MN821 N$6838 N$6836 GND GND n L=2u W=3u
        MP825 N$6836 N$6931 N$6835 VDD p L=2u W=3u
        MP824 N$6836 N$6823 N$6834 VDD p L=2u W=3u
        MP823 N$6835 N$6890 N$6834 VDD p L=2u W=3u
        MP822 N$6834 N$6890 VDD VDD p L=2u W=3u
        MP821 N$6834 N$6931 VDD VDD p L=2u W=3u
        MN820 OUT5 N$6829 GND GND n L=2u W=3u
        MP571 N$6469 N$6471 N$6467 VDD p L=2u W=6u
        MN571 N$6467 CK N$6469 GND n L=2u W=6u
        MN570 N$6469 N$6468 GND GND n L=2u W=6u
        MP570 N$6469 N$6468 VDD VDD p L=2u W=6u
        MN816 N$6831 N$6925 N$6832 GND n L=2u W=3u
        MN815 N$6830 N$6808 GND GND n L=2u W=3u
        MN814 N$6830 N$6867 GND GND n L=2u W=3u
        MN813 N$6830 N$6925 GND GND n L=2u W=3u
        MP574 N$6465 N$6467 VDD VDD p L=2u W=6u
        MN573 N$6910 N$6465 GND GND n L=2u W=6u
        MP573 N$6910 N$6465 VDD VDD p L=2u W=6u
        MP816 N$6827 N$6925 N$6826 VDD p L=2u W=3u
        MN512 N$6779 N$6887 GND GND n L=2u W=3u
        MN511 N$6780 N$6887 GND GND n L=2u W=3u
        MP813 N$6826 N$6808 VDD VDD p L=2u W=3u
        MP812 N$6823 N$6821 VDD VDD p L=2u W=3u
        MN812 N$6821 N$6925 N$6825 GND n L=2u W=3u
        MN811 N$6824 N$6867 GND GND n L=2u W=3u
        MN810 N$6825 N$6867 GND GND n L=2u W=3u
        MN809 N$6821 N$6808 N$6824 GND n L=2u W=3u
        MN808 N$6824 N$6925 GND GND n L=2u W=3u
        MN807 N$6823 N$6821 GND GND n L=2u W=3u
        MP811 N$6821 N$6925 N$6820 VDD p L=2u W=3u
        MP810 N$6821 N$6808 N$6819 VDD p L=2u W=3u
        MP809 N$6820 N$6867 N$6819 VDD p L=2u W=3u
        MP808 N$6819 N$6867 VDD VDD p L=2u W=3u
        MP807 N$6819 N$6925 VDD VDD p L=2u W=3u
        MN806 OUT4 N$6814 GND GND n L=2u W=3u
        MP806 OUT4 N$6814 VDD VDD p L=2u W=3u
        MN805 N$6814 N$6793 N$6816 GND n L=2u W=3u
        MN834 OUT6 N$6844 GND GND n L=2u W=3u
        MP834 OUT6 N$6844 VDD VDD p L=2u W=3u
        MN833 N$6844 N$6823 N$6846 GND n L=2u W=3u
        MN800 N$6815 N$6889 GND GND n L=2u W=3u
        MN799 N$6815 N$6924 GND GND n L=2u W=3u
        MP805 N$6814 N$6806 N$6811 VDD p L=2u W=3u
        MP804 N$6814 N$6793 N$6813 VDD p L=2u W=3u
        MN828 N$6845 N$6890 GND GND n L=2u W=3u
        MN827 N$6845 N$6931 GND GND n L=2u W=3u
        MP833 N$6844 N$6836 N$6841 VDD p L=2u W=3u
        MP800 N$6811 N$6924 VDD VDD p L=2u W=3u
        MN380 N$6750 N$6221 GND GND n L=2u W=3u
        MN379 N$6749 N$6747 GND GND n L=2u W=3u
        MN783 N$6794 N$6888 GND GND n L=2u W=3u
        MN782 N$6795 N$6888 GND GND n L=2u W=3u
        MN781 N$6791 N$6865 N$6794 GND n L=2u W=3u
        MN780 N$6794 N$6923 GND GND n L=2u W=3u
        MN779 N$6793 N$6791 GND GND n L=2u W=3u
        MP783 N$6791 N$6923 N$6790 VDD p L=2u W=3u
        MP782 N$6791 N$6865 N$6789 VDD p L=2u W=3u
        MP781 N$6790 N$6888 N$6789 VDD p L=2u W=3u
        MP780 N$6789 N$6888 VDD VDD p L=2u W=3u
        MP779 N$6789 N$6923 VDD VDD p L=2u W=3u
        MN778 OUT2 N$6784 GND GND n L=2u W=3u
        MP778 OUT2 N$6784 VDD VDD p L=2u W=3u
        MN777 N$6784 N$6764 N$6786 GND n L=2u W=3u
        MN776 N$6784 N$6777 N$6785 GND n L=2u W=3u
        MN775 N$6787 N$6887 GND GND n L=2u W=3u
        MN774 N$6786 N$6922 N$6787 GND n L=2u W=3u
        MP820 OUT5 N$6829 VDD VDD p L=2u W=3u
        MN819 N$6829 N$6808 N$6831 GND n L=2u W=3u
        MN818 N$6829 N$6821 N$6830 GND n L=2u W=3u
        MN817 N$6832 N$6867 GND GND n L=2u W=3u
        MP776 N$6784 N$6764 N$6783 VDD p L=2u W=3u
        MP775 N$6783 N$6887 N$6782 VDD p L=2u W=3u
        MP774 N$6782 N$6922 N$6781 VDD p L=2u W=3u
        MP516 N$6781 N$6887 VDD VDD p L=2u W=3u
        MP819 N$6829 N$6821 N$6826 VDD p L=2u W=3u
        MP818 N$6829 N$6808 N$6828 VDD p L=2u W=3u
        MP817 N$6828 N$6867 N$6827 VDD p L=2u W=3u
        MN513 N$6777 N$6922 N$6780 GND n L=2u W=3u
        MN46 N$1718 GND GND GND n L=2u W=3u
        MN45 N$1715 N$1699 N$1717 GND n L=2u W=3u
        MN394 N$6765 N$6921 GND GND n L=2u W=3u
        MN393 N$6764 N$6762 GND GND n L=2u W=3u
        MP397 N$6762 N$6921 N$6761 VDD p L=2u W=3u
        MP396 N$6762 N$6749 N$6760 VDD p L=2u W=3u
        MP395 N$6761 N$6696 N$6760 VDD p L=2u W=3u
        MP394 N$6760 N$6696 VDD VDD p L=2u W=3u
        MP393 N$6760 N$6921 VDD VDD p L=2u W=3u
        MN392 OUT0 N$6755 GND GND n L=2u W=3u
        MP392 OUT0 N$6755 VDD VDD p L=2u W=3u
        MN391 N$6755 GND N$6757 GND n L=2u W=3u
        MN390 N$6755 N$6747 N$6756 GND n L=2u W=3u
        MN389 N$6758 N$6900 GND GND n L=2u W=3u
        MN388 N$6757 N$6221 N$6758 GND n L=2u W=3u
        MN387 N$6756 GND GND GND n L=2u W=3u
        MN386 N$6756 N$6900 GND GND n L=2u W=3u
        MN385 N$6756 N$6221 GND GND n L=2u W=3u
        MN804 N$6814 N$6806 N$6815 GND n L=2u W=3u
        MN803 N$6817 N$6889 GND GND n L=2u W=3u
        MN802 N$6816 N$6924 N$6817 GND n L=2u W=3u
        MN801 N$6815 N$6793 GND GND n L=2u W=3u
        MP387 N$6752 N$6900 VDD VDD p L=2u W=3u
        MP386 N$6752 N$6221 VDD VDD p L=2u W=3u
        MP385 N$6752 GND VDD VDD p L=2u W=3u
        MP384 N$6749 N$6747 VDD VDD p L=2u W=3u
        MP803 N$6813 N$6889 N$6812 VDD p L=2u W=3u
        MP802 N$6812 N$6924 N$6811 VDD p L=2u W=3u
        MP801 N$6811 N$6889 VDD VDD p L=2u W=3u
        MN381 N$6747 GND N$6750 GND n L=2u W=3u
        MP357 N$6248 N$6689 N$6234 VDD p L=2u W=5u
        MN356 N$6234 N$6689 GND GND n L=2u W=5u
        MN44 N$1717 N$6243 GND GND n L=2u W=3u
        MN355 N$6266 N$6689 GND GND n L=2u W=5u
        MP355 N$6266 N$6689 VDD VDD p L=2u W=5u
        MN354 N$6235 N$6266 N$6246 GND n L=2u W=5u
        MP358 GND N$6266 N$6233 VDD p L=2u W=5u
        MN358 N$6233 N$6689 GND GND n L=2u W=5u
        MP359 N$6250 N$6689 N$6233 VDD p L=2u W=5u
        MN359 N$6233 N$6266 N$6250 GND n L=2u W=5u
        MP353 GND N$6266 N$6235 VDD p L=2u W=5u
        MP158 N$6218 N$6217 N$6214 VDD p L=2u W=6u
        MN158 N$6214 CK N$6218 GND n L=2u W=6u
        MP157 N$5078 CK N$6218 VDD p L=2u W=6u
        MN157 N$6218 N$6217 N$5078 GND n L=2u W=6u
        MN406 N$6619 N$6622 GND GND n L=2u W=3u
        MN134 N$5049 N$6651 N$3358 GND n L=2u W=5u
        MP62 N$1734 N$1732 VDD VDD p L=2u W=3u
        MP64 N$1737 N$6236 VDD VDD p L=2u W=3u
        MP391 N$6755 N$6747 N$6752 VDD p L=2u W=3u
        MP390 N$6755 GND N$6754 VDD p L=2u W=3u
        MP389 N$6754 N$6900 N$6753 VDD p L=2u W=3u
        MP388 N$6753 N$6221 N$6752 VDD p L=2u W=3u
        MN243 N$6223 N$6232 GND GND n L=2u W=6u
        MN244 N$4416 N$5896 N$4418 GND n L=2u W=6u
        MN133 N$5049 N$6933 N$1726 GND n L=2u W=5u
        MN384 N$6747 N$6221 N$6751 GND n L=2u W=3u
        MN383 N$6750 N$6900 GND GND n L=2u W=3u
        MN382 N$6751 N$6900 GND GND n L=2u W=3u
        MN93 N$1777 N$1752 GND GND n L=2u W=3u
        MP246 N$6270 N$6232 N$4413 VDD p L=2u W=6u
        MN246 N$4413 N$5896 N$6270 GND n L=2u W=6u
        MP71 N$1746 N$6255 VDD VDD p L=2u W=3u
        MN245 N$4416 N$6232 GND GND n L=2u W=6u
        MP244 N$4418 N$6232 N$4416 VDD p L=2u W=6u
        MP408 N$6623 N$6624 N$6626 VDD p L=2u W=3u
        MP407 N$6626 N$6624 VDD VDD p L=2u W=3u
        MP406 N$6626 N$6625 VDD VDD p L=2u W=3u
        MP409 N$6622 N$6621 N$6626 VDD p L=2u W=3u
        MN146 N$5065 N$6651 N$6634 GND n L=2u W=5u
        MN20 N$1274 N$6234 N$1278 GND n L=2u W=3u
        MN55 N$1722 N$1699 N$1724 GND n L=2u W=3u
        MP13 N$855 N$245 N$231 VDD p L=2u W=3u
        MN8 N$239 GND GND GND n L=2u W=3u
        MP57 N$1728 N$6236 VDD VDD p L=2u W=3u
        MN25 N$1285 GND GND GND n L=2u W=3u
        MN24 N$1284 N$6234 N$1285 GND n L=2u W=3u
        MN23 N$1283 N$5 GND GND n L=2u W=3u
        MN22 N$1283 GND GND GND n L=2u W=3u
        MP79 N$1755 N$6223 VDD VDD p L=2u W=3u
        MN41 N$1705 N$1276 N$1707 GND n L=2u W=3u
        MN38 N$1707 N$6233 N$1708 GND n L=2u W=3u
        MN139 N$5057 N$6933 N$1762 GND n L=2u W=5u
        MN36 N$1706 GND GND GND n L=2u W=3u
        MN360 N$6243 N$6689 GND GND n L=2u W=5u
        MP360 GND N$6266 N$6243 VDD p L=2u W=5u
        MP21 N$1279 N$5 VDD VDD p L=2u W=3u
        MP20 N$1276 N$1274 VDD VDD p L=2u W=3u
        MN71 N$1752 N$1750 GND GND n L=2u W=3u
        MP75 N$1750 N$6255 N$1749 VDD p L=2u W=3u
        MP410 N$6622 N$6625 N$6623 VDD p L=2u W=3u
        MN97 N$1776 N$1752 N$1778 GND n L=2u W=3u
        MP107 N$1791 N$4416 VDD VDD p L=2u W=3u
        MP106 N$1791 N$6244 VDD VDD p L=2u W=3u
        MP165 N$6217 CK VDD VDD p L=2u W=5u
        MN17 N$1274 N$5 N$1277 GND n L=2u W=3u
        MN18 N$1278 GND GND GND n L=2u W=3u
        MP23 N$1279 GND VDD VDD p L=2u W=3u
        MN13 N$855 GND N$241 GND n L=2u W=3u
        MP42 N$1709 N$1705 VDD VDD p L=2u W=3u
        MN98 N$1780 N$1776 GND GND n L=2u W=3u
        MP70 N$3358 N$1740 VDD VDD p L=2u W=3u
        MN50 N$1723 GND GND GND n L=2u W=3u
        MN96 N$1776 N$1768 N$1777 GND n L=2u W=3u
        MN95 N$1779 N$4413 GND GND n L=2u W=3u
        MP39 N$1704 GND N$1703 VDD p L=2u W=3u
        MN68 N$1740 N$1732 N$1741 GND n L=2u W=3u
        MN67 N$1743 N$6225 GND GND n L=2u W=3u
        MN66 N$1742 N$6236 N$1743 GND n L=2u W=3u
        MP95 N$1775 N$4413 N$1774 VDD p L=2u W=3u
        MP96 N$1776 N$1752 N$1775 VDD p L=2u W=3u
        MP97 N$1776 N$1768 N$1773 VDD p L=2u W=3u
        MP90 N$1770 N$1768 VDD VDD p L=2u W=3u
        MN88 N$1772 N$4413 GND GND n L=2u W=3u
        MN89 N$1771 N$4413 GND GND n L=2u W=3u
        MN58 N$1735 N$6236 GND GND n L=2u W=3u
        MP93 N$1773 N$4413 VDD VDD p L=2u W=3u
        MP94 N$1774 N$6238 N$1773 VDD p L=2u W=3u
        MN49 N$1723 N$6243 GND GND n L=2u W=3u
        MP368 GND N$6266 N$6244 VDD p L=2u W=5u
        MN367 N$6238 N$6266 N$6259 GND n L=2u W=5u
        MP367 N$6259 N$6689 N$6238 VDD p L=2u W=5u
        MP52 N$1720 N$6243 N$1719 VDD p L=2u W=3u
        MN33 N$1700 GND GND GND n L=2u W=3u
        MP34 N$1699 N$1697 VDD VDD p L=2u W=3u
        MN81 N$1761 N$6223 GND GND n L=2u W=3u
        MN104 N$1786 N$6244 N$1790 GND n L=2u W=3u
        MN103 N$1789 N$4416 GND GND n L=2u W=3u
        MN102 N$1790 N$4416 GND GND n L=2u W=3u
        MP2 N$209 GND VDD VDD p L=2u W=3u
        MP25 N$1281 GND N$1280 VDD p L=2u W=3u
        MP26 N$1282 N$5 N$1281 VDD p L=2u W=3u
        MN109 N$1797 N$4416 GND GND n L=2u W=3u
        MN108 N$1796 N$6244 N$1797 GND n L=2u W=3u
        MN73 N$1750 N$1734 N$1753 GND n L=2u W=3u
        MP48 N$1489 N$1715 VDD VDD p L=2u W=3u
        MP49 N$1719 N$1699 VDD VDD p L=2u W=3u
        MP50 N$1719 N$6243 VDD VDD p L=2u W=3u
        MP51 N$1719 GND VDD VDD p L=2u W=3u
        MP38 N$1703 N$6233 N$1702 VDD p L=2u W=3u
        MN11 N$236 GND GND GND n L=2u W=3u
        MN1 N$5 N$245 GND GND n L=2u W=3u
        MP6 N$5 N$245 VDD VDD p L=2u W=3u
        MP46 N$1715 N$1699 N$1711 VDD p L=2u W=3u
        MN69 N$1740 N$1489 N$1742 GND n L=2u W=3u
        MN105 N$1795 N$6244 GND GND n L=2u W=3u
        MP161 N$6214 N$6217 N$6212 VDD p L=2u W=6u
        MN161 N$6212 CK N$6214 GND n L=2u W=6u
        MN160 N$6214 N$6213 GND GND n L=2u W=6u
        MP108 N$1792 N$6244 N$1791 VDD p L=2u W=3u
        MP133 N$1726 N$6651 N$5049 VDD p L=2u W=5u
        MN131 N$5045 N$6651 N$1726 GND n L=2u W=5u
        MP105 N$1791 N$1770 VDD VDD p L=2u W=3u
        MN94 N$1778 N$6238 N$1779 GND n L=2u W=3u
        MN80 N$1760 N$6255 N$1761 GND n L=2u W=3u
        MN79 N$1759 N$1734 GND GND n L=2u W=3u
        MN78 N$1759 N$6223 GND GND n L=2u W=3u
        MN77 N$1759 N$6255 GND GND n L=2u W=3u
        MP83 N$1758 N$1750 N$1755 VDD p L=2u W=3u
        MP18 N$1274 N$5 N$1270 VDD p L=2u W=3u
        MP41 N$1705 N$1697 N$1702 VDD p L=2u W=3u
        MN48 N$1715 N$6243 N$1718 GND n L=2u W=3u
        MN57 N$1734 N$1732 GND GND n L=2u W=3u
        MN112 N$1798 N$1794 GND GND n L=2u W=3u
        MP112 N$1798 N$1794 VDD VDD p L=2u W=3u
        MN111 N$1794 N$1770 N$1796 GND n L=2u W=3u
        MN110 N$1794 N$1786 N$1795 GND n L=2u W=3u
        MP15 N$1270 N$6234 VDD VDD p L=2u W=3u
        MN91 N$1777 N$6238 GND GND n L=2u W=3u
        MP24 N$1280 N$6234 N$1279 VDD p L=2u W=3u
        MN74 N$1754 N$6223 GND GND n L=2u W=3u
        MN59 N$1732 N$1489 N$1735 GND n L=2u W=3u
        MP19 N$1274 N$6234 N$1273 VDD p L=2u W=3u
        MN31 N$1697 N$1276 N$1700 GND n L=2u W=3u
        MN30 N$1700 N$6233 GND GND n L=2u W=3u
        MP17 N$1273 GND N$1270 VDD p L=2u W=3u
        MP55 N$1722 N$1715 N$1719 VDD p L=2u W=3u
        MP54 N$1722 N$1699 N$1721 VDD p L=2u W=3u
        MP53 N$1721 GND N$1720 VDD p L=2u W=3u
        MN32 N$1701 GND GND GND n L=2u W=3u
        MN766 N$6958 N$6691 GND GND n L=2u W=5u
        MN747 N$6958 N$6690 GND GND n L=2u W=5u
        MN198 N$6277 N$6286 GND GND n L=2u W=3u
        MN745 N$6958 N$6685 GND GND n L=2u W=5u
        MN744 N$6958 N$6689 GND GND n L=2u W=5u
        MP766 N$6958 N$6691 N$6303 VDD p L=2u W=5u
        MP173 N$6297 N$6301 VDD VDD p L=2u W=6u
        MP172 N$6301 N$6300 N$6298 VDD p L=2u W=6u
        MN172 N$6298 CK N$6301 GND n L=2u W=6u
        MP171 N$6299 CK N$6301 VDD p L=2u W=6u
        MN171 N$6301 N$6300 N$6299 GND n L=2u W=6u
        MN767 N$8380 N$6958 GND GND n L=2u W=5u
        MP176 N$6296 CK N$6494 VDD p L=2u W=6u
        MN176 N$6494 N$6300 N$6296 GND n L=2u W=6u
        MP175 N$6298 N$6300 N$6296 VDD p L=2u W=6u
        MN175 N$6296 CK N$6298 GND n L=2u W=6u
        MN174 N$6298 N$6297 GND GND n L=2u W=6u
        MP174 N$6298 N$6297 VDD VDD p L=2u W=6u
        MN173 N$6297 N$6301 GND GND n L=2u W=6u
        MN179 N$6300 CK GND GND n L=2u W=5u
        MP771 N$6286 H0 VDD VDD p L=2u W=3u
        MP473 N$6553 N$6558 VDD VDD p L=2u W=5u
        MN473 N$6550 N$6558 GND GND n L=2u W=5u
        MN773 N$6572 N$6497 N$6519 GND n L=2u W=5u
        MN177 N$6494 N$6295 GND GND n L=2u W=6u
        MP177 N$6494 N$6295 VDD VDD p L=2u W=6u
        MN182 N$6291 N$6294 GND GND n L=2u W=6u
        MP182 N$6291 N$6294 VDD VDD p L=2u W=6u
        MN16 N$1277 N$6234 GND GND n L=2u W=3u
        MP33 N$1697 N$6233 N$1696 VDD p L=2u W=3u
        MP32 N$1697 N$1276 N$1693 VDD p L=2u W=3u
        MN180 N$6294 N$6293 N$6545 GND n L=2u W=6u
        MN754 N$6689 N$6313 GND GND n L=2u W=6u
        MP754 N$6689 N$6313 VDD VDD p L=2u W=6u
        MP184 N$6292 N$6293 N$6290 VDD p L=2u W=6u
        MN753 N$6689 N$6317 N$6314 GND n L=2u W=6u
        MP752 N$6316 N$6317 N$6314 VDD p L=2u W=6u
        MN752 N$6314 CK N$6316 GND n L=2u W=6u
        MP757 N$6328 CK N$6312 VDD p L=2u W=6u
        MN757 N$6312 N$6311 N$6328 GND n L=2u W=6u
        MN756 N$6317 CK GND GND n L=2u W=5u
        MP756 N$6317 CK VDD VDD p L=2u W=5u
        MN755 N$6313 N$6314 GND GND n L=2u W=6u
        MP761 N$6310 N$6311 N$6308 VDD p L=2u W=6u
        MN761 N$6308 CK N$6310 GND n L=2u W=6u
        MN760 N$6310 N$6309 GND GND n L=2u W=6u
        MP760 N$6310 N$6309 VDD VDD p L=2u W=6u
        MN759 N$6309 N$6312 GND GND n L=2u W=6u
        MP759 N$6309 N$6312 VDD VDD p L=2u W=6u
        MP758 N$6312 N$6311 N$6310 VDD p L=2u W=6u
        MN758 N$6310 CK N$6312 GND n L=2u W=6u
        MP764 N$6692 N$6308 VDD VDD p L=2u W=6u
        MN194 N$6282 N$6286 GND GND n L=2u W=3u
        MN193 N$6284 C0 N$6283 GND n L=2u W=3u
        MN192 N$6283 N$6542 GND GND n L=2u W=3u
        MN191 N$6621 N$6284 GND GND n L=2u W=3u
        MP747 N$6303 N$6690 N$6304 VDD p L=2u W=5u
        MP746 N$6304 N$6328 N$6305 VDD p L=2u W=5u
        MP745 N$6305 N$6685 N$6306 VDD p L=2u W=5u
        MP744 N$6306 N$6689 VDD VDD p L=2u W=5u
        MP198 N$6281 N$6542 VDD VDD p L=2u W=3u
        MP197 N$6281 C0 VDD VDD p L=2u W=3u
        MP196 N$6621 N$6284 VDD VDD p L=2u W=3u
        MP767 N$8380 N$6958 VDD VDD p L=2u W=5u
        MP734 N$6332 CK VDD VDD p L=2u W=5u
        MN733 N$6688 N$6329 GND GND n L=2u W=6u
        MN746 N$6958 N$6328 GND GND n L=2u W=5u
        MP733 N$6688 N$6329 VDD VDD p L=2u W=6u
        MN732 N$6328 N$6688 GND GND n L=2u W=6u
        MN738 N$6323 N$6322 GND GND n L=2u W=6u
        MP738 N$6323 N$6322 VDD VDD p L=2u W=6u
        MN737 N$6322 N$6326 GND GND n L=2u W=6u
        MP737 N$6322 N$6326 VDD VDD p L=2u W=6u
        MP736 N$6326 N$6325 N$6323 VDD p L=2u W=6u
        MN736 N$6323 CK N$6326 GND n L=2u W=6u
        MP735 N$6690 CK N$6326 VDD p L=2u W=6u
        MN741 N$6691 N$6319 GND GND n L=2u W=6u
        MP741 N$6691 N$6319 VDD VDD p L=2u W=6u
        MP740 N$6321 CK N$6691 VDD p L=2u W=6u
        MN740 N$6691 N$6325 N$6321 GND n L=2u W=6u
        MP739 N$6323 N$6325 N$6321 VDD p L=2u W=6u
        MN739 N$6321 CK N$6323 GND n L=2u W=6u
        MP748 N$6682 CK N$6318 VDD p L=2u W=6u
        MN748 N$6318 N$6317 N$6682 GND n L=2u W=6u
        MP179 N$6300 CK VDD VDD p L=2u W=5u
        MN178 N$6295 N$6296 GND GND n L=2u W=6u
        MP178 N$6295 N$6296 VDD VDD p L=2u W=6u
        MP742 N$6319 N$6321 VDD VDD p L=2u W=6u
        MN751 N$6316 N$6315 GND GND n L=2u W=6u
        MP751 N$6316 N$6315 VDD VDD p L=2u W=6u
        MN750 N$6315 N$6318 GND GND n L=2u W=6u
        MP181 N$6294 N$6293 N$6292 VDD p L=2u W=6u
        MN181 N$6292 CK N$6294 GND n L=2u W=6u
        MP180 N$6545 CK N$6294 VDD p L=2u W=6u
        MP755 N$6313 N$6314 VDD VDD p L=2u W=6u
        MP718 N$6341 N$6340 N$6338 VDD p L=2u W=6u
        MN718 N$6338 CK N$6341 GND n L=2u W=6u
        MP753 N$6314 CK N$6689 VDD p L=2u W=6u
        MN717 N$6341 N$6340 N$6689 GND n L=2u W=6u
        MN716 N$6347 CK GND GND n L=2u W=5u
        MP722 N$6336 CK N$6685 VDD p L=2u W=6u
        MN722 N$6685 N$6340 N$6336 GND n L=2u W=6u
        MP721 N$6338 N$6340 N$6336 VDD p L=2u W=6u
        MN721 N$6336 CK N$6338 GND n L=2u W=6u
        MN720 N$6338 N$6337 GND GND n L=2u W=6u
        MP720 N$6338 N$6337 VDD VDD p L=2u W=6u
        MN725 N$6340 CK GND GND n L=2u W=5u
        MP725 N$6340 CK VDD VDD p L=2u W=5u
        MN724 N$6687 N$6336 GND GND n L=2u W=6u
        MP724 N$6687 N$6336 VDD VDD p L=2u W=6u
        MN723 N$6685 N$6687 GND GND n L=2u W=6u
        MP723 N$6685 N$6687 VDD VDD p L=2u W=6u
        MN728 N$6330 N$6333 GND GND n L=2u W=6u
        MP728 N$6330 N$6333 VDD VDD p L=2u W=6u
        MP727 N$6333 N$6332 N$6331 VDD p L=2u W=6u
        MN763 N$6690 N$6692 GND GND n L=2u W=6u
        MP763 N$6690 N$6692 VDD VDD p L=2u W=6u
        MP762 N$6308 CK N$6690 VDD p L=2u W=6u
        MN762 N$6690 N$6311 N$6308 GND n L=2u W=6u
        MP731 N$6329 CK N$6328 VDD p L=2u W=6u
        MN731 N$6328 N$6332 N$6329 GND n L=2u W=6u
        MP730 N$6331 N$6332 N$6329 VDD p L=2u W=6u
        MN730 N$6329 CK N$6331 GND n L=2u W=6u
        MN765 N$6311 CK GND GND n L=2u W=5u
        MP765 N$6311 CK VDD VDD p L=2u W=5u
        MN764 N$6692 N$6308 GND GND n L=2u W=6u
        MN734 N$6332 CK GND GND n L=2u W=5u
        MN702 N$6352 N$6351 GND GND n L=2u W=6u
        MP702 N$6352 N$6351 VDD VDD p L=2u W=6u
        MP701 N$6351 N$6354 VDD VDD p L=2u W=6u
        MN706 N$6349 N$6350 GND GND n L=2u W=6u
        MP706 N$6349 N$6350 VDD VDD p L=2u W=6u
        MN705 N$6270 N$6349 GND GND n L=2u W=6u
        MP705 N$6270 N$6349 VDD VDD p L=2u W=6u
        MP704 N$6350 CK N$6270 VDD p L=2u W=6u
        MN704 N$6270 N$6353 N$6350 GND n L=2u W=6u
        MP710 N$6345 N$6348 VDD VDD p L=2u W=6u
        MP709 N$6348 N$6347 N$6346 VDD p L=2u W=6u
        MN709 N$6346 CK N$6348 GND n L=2u W=6u
        MP708 N$6368 CK N$6348 VDD p L=2u W=6u
        MN708 N$6348 N$6347 N$6368 GND n L=2u W=6u
        MN707 N$6353 CK GND GND n L=2u W=5u
        MP707 N$6353 CK VDD VDD p L=2u W=5u
        MN713 N$4418 N$6347 N$6344 GND n L=2u W=6u
        MP712 N$6346 N$6347 N$6344 VDD p L=2u W=6u
        MN712 N$6344 CK N$6346 GND n L=2u W=6u
        MN743 N$6325 CK GND GND n L=2u W=5u
        MP743 N$6325 CK VDD VDD p L=2u W=5u
        MN742 N$6319 N$6321 GND GND n L=2u W=6u
        MP716 N$6347 CK VDD VDD p L=2u W=5u
        MN715 N$6343 N$6344 GND GND n L=2u W=6u
        MP715 N$6343 N$6344 VDD VDD p L=2u W=6u
        MN714 N$4418 N$6343 GND GND n L=2u W=6u
        MP750 N$6315 N$6318 VDD VDD p L=2u W=6u
        MP749 N$6318 N$6317 N$6316 VDD p L=2u W=6u
        MN749 N$6316 CK N$6318 GND n L=2u W=6u
        MP719 N$6337 N$6341 VDD VDD p L=2u W=6u
        MN686 N$6268 N$9223 N$6362 GND n L=2u W=6u
        MP685 N$6364 N$9223 N$6362 VDD p L=2u W=6u
        MP717 N$6689 CK N$6341 VDD p L=2u W=6u
        MP690 N$6370 CK N$6360 VDD p L=2u W=6u
        MN690 N$6360 N$6359 N$6370 GND n L=2u W=6u
        MN689 N$9223 CK GND GND n L=2u W=5u
        MP689 N$9223 CK VDD VDD p L=2u W=5u
        MN688 N$6361 N$6362 GND GND n L=2u W=6u
        MP688 N$6361 N$6362 VDD VDD p L=2u W=6u
        MN694 N$6356 CK N$6358 GND n L=2u W=6u
        MN693 N$6358 N$6357 GND GND n L=2u W=6u
        MP693 N$6358 N$6357 VDD VDD p L=2u W=6u
        MN692 N$6357 N$6360 GND GND n L=2u W=6u
        MP692 N$6357 N$6360 VDD VDD p L=2u W=6u
        MP691 N$6360 N$6359 N$6358 VDD p L=2u W=6u
        MN691 N$6358 CK N$6360 GND n L=2u W=6u
        MP697 N$6355 N$6356 VDD VDD p L=2u W=6u
        MN696 N$6269 N$6355 GND GND n L=2u W=6u
        MP696 N$6269 N$6355 VDD VDD p L=2u W=6u
        MN727 N$6331 CK N$6333 GND n L=2u W=6u
        MP726 N$6685 CK N$6333 VDD p L=2u W=6u
        MN726 N$6333 N$6332 N$6685 GND n L=2u W=6u
        MP732 N$6328 N$6688 VDD VDD p L=2u W=6u
        MN700 N$6352 CK N$6354 GND n L=2u W=6u
        MP699 N$6369 CK N$6354 VDD p L=2u W=6u
        MN699 N$6354 N$6353 N$6369 GND n L=2u W=6u
        MN698 N$6359 CK GND GND n L=2u W=5u
        MN729 N$6331 N$6330 GND GND n L=2u W=6u
        MP729 N$6331 N$6330 VDD VDD p L=2u W=6u
        MN735 N$6326 N$6325 N$6690 GND n L=2u W=6u
        MN703 N$6350 CK N$6352 GND n L=2u W=6u
        MP644 N$6393 N$6397 VDD VDD p L=2u W=3u
        MN643 N$6397 N$6418 N$6395 GND n L=2u W=3u
        MP675 N$6408 N$6376 N$6370 VDD p L=2u W=5u
        MN641 N$6394 N$6406 GND GND n L=2u W=3u
        MN640 N$6395 H2 N$6394 GND n L=2u W=3u
        MN639 N$6396 N$6418 GND GND n L=2u W=3u
        MN645 COUTHK-SK N$6389 GND GND n L=2u W=3u
        MP649 N$6389 H3 N$6390 VDD p L=2u W=3u
        MP648 N$6389 N$6403 N$6392 VDD p L=2u W=3u
        MP647 N$6390 N$6391 N$6392 VDD p L=2u W=3u
        MP646 N$6392 N$6391 VDD VDD p L=2u W=3u
        MP645 N$6392 H3 VDD VDD p L=2u W=3u
        MP650 COUTHK-SK N$6389 VDD VDD p L=2u W=3u
        MN650 N$6389 H3 N$6386 GND n L=2u W=3u
        MN649 N$6387 N$6391 GND GND n L=2u W=3u
        MN648 N$6386 N$6391 GND GND n L=2u W=3u
        MN647 N$6389 N$6403 N$6387 GND n L=2u W=3u
        MN646 N$6387 H3 GND GND n L=2u W=3u
        MP657 N$6382 N$6389 N$6385 VDD p L=2u W=3u
        MP656 N$6382 N$6403 N$6383 VDD p L=2u W=3u
        MN711 N$6346 N$6345 GND GND n L=2u W=6u
        MP711 N$6346 N$6345 VDD VDD p L=2u W=6u
        MN710 N$6345 N$6348 GND GND n L=2u W=6u
        MP684 N$6364 N$6363 VDD VDD p L=2u W=6u
        MN683 N$6363 N$6366 GND GND n L=2u W=6u
        MP683 N$6363 N$6366 VDD VDD p L=2u W=6u
        MP682 N$6366 N$9223 N$6364 VDD p L=2u W=6u
        MP714 N$4418 N$6343 VDD VDD p L=2u W=6u
        MP713 N$6344 CK N$4418 VDD p L=2u W=6u
        MN719 N$6337 N$6341 GND GND n L=2u W=6u
        MP686 N$6362 CK N$6268 VDD p L=2u W=6u
        MN626 N$6410 H1 N$6409 GND n L=2u W=3u
        MN625 N$6411 N$8383 GND GND n L=2u W=3u
        MN658 N$6378 N$6382 GND GND n L=2u W=3u
        MN623 N$6411 H1 GND GND n L=2u W=3u
        MP629 N$6412 N$6419 N$6415 VDD p L=2u W=3u
        MP632 N$6407 N$6406 VDD VDD p L=2u W=3u
        MP631 N$6407 H2 VDD VDD p L=2u W=3u
        MN630 N$6408 N$6412 GND GND n L=2u W=3u
        MP630 N$6408 N$6412 VDD VDD p L=2u W=3u
        MN629 N$6412 N$8383 N$6410 GND n L=2u W=3u
        MN628 N$6412 N$6419 N$6411 GND n L=2u W=3u
        MN633 N$6404 N$6418 N$6402 GND n L=2u W=3u
        MN632 N$6402 H2 GND GND n L=2u W=3u
        MN631 N$6403 N$6404 GND GND n L=2u W=3u
        MP635 N$6404 H2 N$6405 VDD p L=2u W=3u
        MP634 N$6404 N$6418 N$6407 VDD p L=2u W=3u
        MP633 N$6405 N$6406 N$6407 VDD p L=2u W=3u
        MP639 N$6400 N$6406 VDD VDD p L=2u W=3u
        MP638 N$6400 H2 VDD VDD p L=2u W=3u
        MN663 N$6479 N$6515 N$9213 GND n L=2u W=5u
        MP669 N$6484 N$6515 N$6462 VDD p L=2u W=5u
        MN668 N$6462 N$6515 N$6443 GND n L=2u W=5u
        MP668 N$6443 N$6376 N$6462 VDD p L=2u W=5u
        MN634 N$6401 N$6406 GND GND n L=2u W=3u
        MN638 N$6396 N$6406 GND GND n L=2u W=3u
        MN637 N$6396 H2 GND GND n L=2u W=3u
        MP643 N$6397 N$6404 N$6400 VDD p L=2u W=3u
        MN671 N$6454 N$6376 N$6483 GND n L=2u W=5u
        MP671 N$6483 N$6515 N$6454 VDD p L=2u W=5u
        MN644 N$6393 N$6397 GND GND n L=2u W=3u
        MP537 N$6658 N$6500 VDD VDD p L=2u W=6u
        MN536 N$9207 N$6658 GND GND n L=2u W=6u
        MP568 N$6472 N$6471 N$6469 VDD p L=2u W=6u
        MP535 N$6500 CK N$9207 VDD p L=2u W=6u
        MN541 N$6542 N$6497 N$6494 GND n L=2u W=5u
        MP541 N$6494 RST N$6542 VDD p L=2u W=5u
        MN540 N$6542 RST A5 GND n L=2u W=5u
        MP540 A5 N$6497 N$6542 VDD p L=2u W=5u
        MN539 N$6499 N$8173 GND GND n L=2u W=6u
        MP539 N$6499 N$8173 VDD VDD p L=2u W=6u
        MN544 N$6625 N$6497 N$6533 GND n L=2u W=5u
        MP544 N$6533 RST N$6625 VDD p L=2u W=5u
        MN543 N$6625 RST GND GND n L=2u W=5u
        MP543 GND N$6497 N$6625 VDD p L=2u W=5u
        MN542 N$6497 RST GND GND n L=2u W=5u
        MP542 N$6497 RST VDD VDD p L=2u W=5u
        MN547 N$6588 RST GND GND n L=2u W=5u
        MP547 GND N$6497 N$6588 VDD p L=2u W=5u
        MN546 N$6605 N$6497 N$6526 GND n L=2u W=5u
        MP655 N$6383 N$6391 N$6384 VDD p L=2u W=3u
        MP654 N$6384 H3 N$6385 VDD p L=2u W=3u
        MP653 N$6385 N$6391 VDD VDD p L=2u W=3u
        MP652 N$6385 H3 VDD VDD p L=2u W=3u
        MP628 N$6412 N$8383 N$6413 VDD p L=2u W=3u
        MP627 N$6413 N$6421 N$6414 VDD p L=2u W=3u
        MP626 N$6414 H1 N$6415 VDD p L=2u W=3u
        MP625 N$6415 N$6421 VDD VDD p L=2u W=3u
        MN653 N$6381 N$6403 GND GND n L=2u W=3u
        MN652 N$6381 N$6391 GND GND n L=2u W=3u
        MN651 N$6381 H3 GND GND n L=2u W=3u
        MN627 N$6409 N$6421 GND GND n L=2u W=3u
        MN521 N$6510 N$6509 N$6550 GND n L=2u W=6u
        MN520 N$6511 N$6516 GND GND n L=2u W=5u
        MN552 N$6485 N$6499 N$6533 GND n L=2u W=5u
        MP520 N$8173 N$6516 VDD VDD p L=2u W=5u
        MP525 N$6508 N$6509 N$6506 VDD p L=2u W=6u
        MN525 N$6506 CK N$6508 GND n L=2u W=6u
        MN524 N$6508 N$6507 GND GND n L=2u W=6u
        MP524 N$6508 N$6507 VDD VDD p L=2u W=6u
        MN523 N$6507 N$6510 GND GND n L=2u W=6u
        MP523 N$6507 N$6510 VDD VDD p L=2u W=6u
        MN528 N$6505 N$6506 GND GND n L=2u W=6u
        MP528 N$6505 N$6506 VDD VDD p L=2u W=6u
        MN527 N$6516 N$6505 GND GND n L=2u W=6u
        MP527 N$6516 N$6505 VDD VDD p L=2u W=6u
        MP526 N$6506 CK N$6516 VDD p L=2u W=6u
        MN526 N$6516 N$6509 N$6506 GND n L=2u W=6u
        MP532 N$6501 N$6504 VDD VDD p L=2u W=6u
        MP531 N$6504 N$6503 N$6502 VDD p L=2u W=6u
        MN531 N$6502 CK N$6504 GND n L=2u W=6u
        MP530 N$6683 CK N$6504 VDD p L=2u W=6u
        MP562 N$6477 N$6480 N$6475 VDD p L=2u W=6u
        MN562 N$6475 CK N$6477 GND n L=2u W=6u
        MN561 N$6477 N$6476 GND GND n L=2u W=6u
        MP561 N$6477 N$6476 VDD VDD p L=2u W=6u
        MP534 N$6502 N$6503 N$6500 VDD p L=2u W=6u
        MN534 N$6500 CK N$6502 GND n L=2u W=6u
        MN533 N$6502 N$6501 GND GND n L=2u W=6u
        MP533 N$6502 N$6501 VDD VDD p L=2u W=6u
        MP565 N$6473 N$6475 VDD VDD p L=2u W=6u
        MN564 HK_SK N$6473 GND GND n L=2u W=6u
        MP564 HK_SK N$6473 VDD VDD p L=2u W=6u
        MN537 N$6658 N$6500 GND GND n L=2u W=6u
        MN479 N$6543 N$6683 N$6625 GND n L=2u W=5u
        MP479 N$6625 N$6548 N$6543 VDD p L=2u W=5u
        MN519 N$8173 N$9207 N$6511 GND n L=2u W=5u
        MN484 N$6536 N$6535 GND GND n L=2u W=6u
        MP484 N$6536 N$6535 VDD VDD p L=2u W=6u
        MN483 N$6535 N$6540 GND GND n L=2u W=6u
        MP483 N$6535 N$6540 VDD VDD p L=2u W=6u
        MP482 N$6540 N$6539 N$6536 VDD p L=2u W=6u
        MN482 N$6536 CK N$6540 GND n L=2u W=6u
        MP488 N$6532 N$6534 VDD VDD p L=2u W=6u
        MN487 N$6533 N$6532 GND GND n L=2u W=6u
        MP487 N$6533 N$6532 VDD VDD p L=2u W=6u
        MP486 N$6534 CK N$6533 VDD p L=2u W=6u
        MN486 N$6533 N$6539 N$6534 GND n L=2u W=6u
        MP485 N$6536 N$6539 N$6534 VDD p L=2u W=6u
        MP491 N$6531 N$6530 N$6529 VDD p L=2u W=6u
        MN491 N$6529 CK N$6531 GND n L=2u W=6u
        MP490 N$6544 CK N$6531 VDD p L=2u W=6u
        MN490 N$6531 N$6530 N$6544 GND n L=2u W=6u
        MN489 N$6539 CK GND GND n L=2u W=5u
        MN530 N$6504 N$6503 N$6683 GND n L=2u W=6u
        MN529 N$6509 CK GND GND n L=2u W=6u
        MP529 N$6509 CK VDD VDD p L=2u W=6u
        MN535 N$9207 N$6503 N$6500 GND n L=2u W=6u
        MN493 N$6529 N$6528 GND GND n L=2u W=6u
        MP493 N$6529 N$6528 VDD VDD p L=2u W=6u
        MN492 N$6528 N$6531 GND GND n L=2u W=6u
        MP492 N$6528 N$6531 VDD VDD p L=2u W=6u
        MN532 N$6501 N$6504 GND GND n L=2u W=6u
        MN538 N$6503 CK GND GND n L=2u W=5u
        MP538 N$6503 CK VDD VDD p L=2u W=5u
        MN496 N$6526 N$6525 GND GND n L=2u W=6u
        MN461 N$6558 N$6562 GND GND n L=2u W=3u
        MN495 N$6526 N$6530 N$6527 GND n L=2u W=6u
        MP467 N$6552 N$6609 N$6555 VDD p L=2u W=6u
        MP466 N$6555 N$6554 N$6553 VDD p L=2u W=6u
        MN465 N$6587 H3 GND GND n L=2u W=3u
        MP465 N$6587 H3 VDD VDD p L=2u W=3u
        MN464 N$6571 GND GND GND n L=2u W=3u
        MN470 N$6547 N$6683 N$6572 GND n L=2u W=5u
        MP470 N$6572 N$6548 N$6547 VDD p L=2u W=5u
        MN469 N$6550 N$6574 GND GND n L=2u W=6u
        MN468 N$6550 N$6591 GND GND n L=2u W=6u
        MN467 N$6550 N$6609 GND GND n L=2u W=6u
        MN466 N$6550 N$6554 GND GND n L=2u W=6u
        MP469 N$6550 N$6574 N$6551 VDD p L=2u W=6u
        MN475 N$6545 N$6683 N$6588 GND n L=2u W=5u
        MP475 N$6588 N$6548 N$6545 VDD p L=2u W=5u
        MN472 N$6548 N$6683 GND GND n L=2u W=5u
        MP472 N$6548 N$6683 VDD VDD p L=2u W=5u
        MP505 N$6519 N$6518 VDD VDD p L=2u W=6u
        MP504 N$6520 CK N$6519 VDD p L=2u W=6u
        MP519 N$8173 N$9207 VDD VDD p L=2u W=5u
        MN518 N$6515 N$6658 GND GND n L=2u W=5u
        MN477 N$6544 N$6683 N$6605 GND n L=2u W=5u
        MP477 N$6605 N$6548 N$6544 VDD p L=2u W=5u
        MN476 N$6545 N$6548 N$6605 GND n L=2u W=5u
        MP476 N$6605 N$6683 N$6545 VDD p L=2u W=5u
        MP522 N$6510 N$6509 N$6508 VDD p L=2u W=6u
        MN522 N$6508 CK N$6510 GND n L=2u W=6u
        MP480 N$6542 N$6683 N$6543 VDD p L=2u W=5u
        MP436 N$6586 N$6587 N$6589 VDD p L=2u W=3u
        MP435 N$6589 N$6587 VDD VDD p L=2u W=3u
        MP468 N$6551 N$6591 N$6552 VDD p L=2u W=6u
        MN433 N$6591 N$6595 GND GND n L=2u W=3u
        MN439 N$6585 N$6588 N$6582 GND n L=2u W=3u
        MN438 N$6583 N$6587 GND GND n L=2u W=3u
        MN437 N$6582 N$6587 GND GND n L=2u W=3u
        MN436 N$6585 N$6601 N$6583 GND n L=2u W=3u
        MN435 N$6583 N$6588 GND GND n L=2u W=3u
        MN434 N$6584 N$6585 GND GND n L=2u W=3u
        MP438 N$6585 N$6588 N$6586 VDD p L=2u W=3u
        MP444 N$6579 N$6587 N$6580 VDD p L=2u W=3u
        MP443 N$6580 N$6588 N$6581 VDD p L=2u W=3u
        MP442 N$6581 N$6587 VDD VDD p L=2u W=3u
        MP441 N$6581 N$6588 VDD VDD p L=2u W=3u
        MP440 N$6581 N$6601 VDD VDD p L=2u W=3u
        MP439 N$6584 N$6585 VDD VDD p L=2u W=3u
        MN444 N$6575 N$6587 GND GND n L=2u W=3u
        MN471 N$6547 N$6548 N$6588 GND n L=2u W=5u
        MP471 N$6588 N$6683 N$6547 VDD p L=2u W=5u
        MN478 N$6544 N$6548 N$6625 GND n L=2u W=5u
        MP478 N$6625 N$6683 N$6544 VDD p L=2u W=5u
        MP446 N$6578 N$6585 N$6581 VDD p L=2u W=3u
        MP445 N$6578 N$6601 N$6579 VDD p L=2u W=3u
        MP449 N$6573 N$6571 VDD VDD p L=2u W=3u
        MP448 N$6573 N$6572 VDD VDD p L=2u W=3u
        MP481 N$6543 CK N$6540 VDD p L=2u W=6u
        MN481 N$6540 N$6539 N$6543 GND n L=2u W=6u
        MN480 N$6543 N$6548 N$6542 GND n L=2u W=5u
        MN445 N$6578 N$6585 N$6577 GND n L=2u W=3u
        MN419 N$6609 N$6613 GND GND n L=2u W=3u
        MN448 N$6683 N$6569 GND GND n L=2u W=3u
        MN418 N$6613 N$6621 N$6611 GND n L=2u W=3u
        MN417 N$6613 N$6622 N$6612 GND n L=2u W=3u
        MN422 N$6602 N$6619 N$6600 GND n L=2u W=3u
        MN421 N$6600 N$6605 GND GND n L=2u W=3u
        MN420 N$6601 N$6602 GND GND n L=2u W=3u
        MP424 N$6602 N$6605 N$6603 VDD p L=2u W=3u
        MP423 N$6602 N$6619 N$6606 VDD p L=2u W=3u
        MP422 N$6603 N$6604 N$6606 VDD p L=2u W=3u
        MP421 N$6606 N$6604 VDD VDD p L=2u W=3u
        MP427 N$6598 N$6605 VDD VDD p L=2u W=3u
        MP426 N$6598 N$6619 VDD VDD p L=2u W=3u
        MP425 N$6601 N$6602 VDD VDD p L=2u W=3u
        MN425 N$6602 N$6605 N$6599 GND n L=2u W=3u
        MN424 N$6600 N$6604 GND GND n L=2u W=3u
        MN423 N$6599 N$6604 GND GND n L=2u W=3u
        MN426 N$6594 N$6605 GND GND n L=2u W=3u
        MP432 N$6595 N$6602 N$6598 VDD p L=2u W=3u
        MP461 N$6558 N$6562 VDD VDD p L=2u W=3u
        MN460 N$6562 N$6584 N$6560 GND n L=2u W=3u
        MN459 N$6562 N$6569 N$6561 GND n L=2u W=3u
        MN458 N$6559 N$6571 GND GND n L=2u W=3u
        MP433 N$6591 N$6595 VDD VDD p L=2u W=3u
        MN432 N$6595 N$6619 N$6593 GND n L=2u W=3u
        MN431 N$6595 N$6602 N$6594 GND n L=2u W=3u
        MN430 N$6592 N$6604 GND GND n L=2u W=3u
        MP463 N$6604 H2 VDD VDD p L=2u W=3u
        MN462 N$6624 H1 GND GND n L=2u W=3u
        MP462 N$6624 H1 VDD VDD p L=2u W=3u
        MP437 N$6585 N$6601 N$6589 VDD p L=2u W=3u
        MP250 N$6203 N$6205 VDD VDD p L=2u W=6u
        MN249 N$6204 N$6203 GND GND n L=2u W=6u
        MP434 N$6589 N$6588 VDD VDD p L=2u W=3u
        MN254 N$6199 N$6202 GND GND n L=2u W=6u
        MP254 N$6199 N$6202 VDD VDD p L=2u W=6u
        MP253 N$6202 N$6201 N$6200 VDD p L=2u W=6u
        MN253 N$6200 CK N$6202 GND n L=2u W=6u
        MP252 N$5045 CK N$6202 VDD p L=2u W=6u
        MN252 N$6202 N$6201 N$5045 GND n L=2u W=6u
        MP258 N$6197 N$6196 VDD VDD p L=2u W=6u
        MP257 N$6198 CK N$6197 VDD p L=2u W=6u
        MN257 N$6197 N$6201 N$6198 GND n L=2u W=6u
        MP256 N$6200 N$6201 N$6198 VDD p L=2u W=6u
        MN256 N$6198 CK N$6200 GND n L=2u W=6u
        MN255 N$6200 N$6199 GND GND n L=2u W=6u
        MP255 N$6200 N$6199 VDD VDD p L=2u W=6u
        MN261 N$6195 N$6194 N$5049 GND n L=2u W=6u
        MP415 N$6615 N$6625 N$6616 VDD p L=2u W=3u
        MP414 N$6616 N$6624 VDD VDD p L=2u W=3u
        MP413 N$6616 N$6625 VDD VDD p L=2u W=3u
        MN443 N$6576 N$6588 N$6575 GND n L=2u W=3u
        MN442 N$6577 N$6601 GND GND n L=2u W=3u
        MN441 N$6577 N$6587 GND GND n L=2u W=3u
        MN440 N$6577 N$6588 GND GND n L=2u W=3u
        MN414 N$6612 N$6621 GND GND n L=2u W=3u
        MN413 N$6612 N$6624 GND GND n L=2u W=3u
        MN412 N$6612 N$6625 GND GND n L=2u W=3u
        MP418 N$6613 N$6622 N$6616 VDD p L=2u W=3u
        MN447 N$6574 N$6578 GND GND n L=2u W=3u
        MP447 N$6574 N$6578 VDD VDD p L=2u W=3u
        MN446 N$6578 N$6601 N$6576 GND n L=2u W=3u
        MN266 N$6190 N$6194 N$6191 GND n L=2u W=6u
        MP265 N$6193 N$6194 N$6191 VDD p L=2u W=6u
        MP419 N$6609 N$6613 VDD VDD p L=2u W=3u
        MP270 N$5053 CK N$6188 VDD p L=2u W=6u
        MN270 N$6188 N$6187 N$5053 GND n L=2u W=6u
        MN269 N$6194 CK GND GND n L=2u W=5u
        MP269 N$6194 CK VDD VDD p L=2u W=5u
        MN268 N$6189 N$6191 GND GND n L=2u W=6u
        MP268 N$6189 N$6191 VDD VDD p L=2u W=6u
        MN273 N$6186 N$6185 GND GND n L=2u W=6u
        MP273 N$6186 N$6185 VDD VDD p L=2u W=6u
        MN272 N$6185 N$6188 GND GND n L=2u W=6u
        MP272 N$6185 N$6188 VDD VDD p L=2u W=6u
        MP271 N$6188 N$6187 N$6186 VDD p L=2u W=6u
        MN271 N$6186 CK N$6188 GND n L=2u W=6u
        MP277 N$6182 N$6184 VDD VDD p L=2u W=6u
        MN276 N$6183 N$6182 GND GND n L=2u W=6u
        MP167 N$6209 N$6208 N$6207 VDD p L=2u W=6u
        MN167 N$6207 CK N$6209 GND n L=2u W=6u
        MP166 N$5073 CK N$6209 VDD p L=2u W=6u
        MP431 N$6595 N$6619 N$6596 VDD p L=2u W=3u
        MP430 N$6596 N$6604 N$6597 VDD p L=2u W=3u
        MP429 N$6597 N$6605 N$6598 VDD p L=2u W=3u
        MP428 N$6598 N$6604 VDD VDD p L=2u W=3u
        MP170 N$6207 N$6208 N$6205 VDD p L=2u W=6u
        MN170 N$6205 CK N$6207 GND n L=2u W=6u
        MN169 N$6207 N$6206 GND GND n L=2u W=6u
        MP169 N$6207 N$6206 VDD VDD p L=2u W=6u
        MN429 N$6593 N$6605 N$6592 GND n L=2u W=3u
        MN428 N$6594 N$6619 GND GND n L=2u W=3u
        MN427 N$6594 N$6604 GND GND n L=2u W=3u
        MN250 N$6203 N$6205 GND GND n L=2u W=6u
        MP282 N$6179 N$6178 VDD VDD p L=2u W=6u
        MN281 N$6178 N$6181 GND GND n L=2u W=6u
        MP249 N$6204 N$6203 VDD VDD p L=2u W=6u
        MN286 N$6175 N$6177 GND GND n L=2u W=6u
        MP286 N$6175 N$6177 VDD VDD p L=2u W=6u
        MN285 N$6176 N$6175 GND GND n L=2u W=6u
        MP285 N$6176 N$6175 VDD VDD p L=2u W=6u
        MP284 N$6177 CK N$6176 VDD p L=2u W=6u
        MN284 N$6176 N$6180 N$6177 GND n L=2u W=6u
        MP290 N$6171 N$6174 VDD VDD p L=2u W=6u
        MP289 N$6174 N$6173 N$6172 VDD p L=2u W=6u
        MN289 N$6172 CK N$6174 GND n L=2u W=6u
        MP288 N$5061 CK N$6174 VDD p L=2u W=6u
        MN288 N$6174 N$6173 N$5061 GND n L=2u W=6u
        MN287 N$6180 CK GND GND n L=2u W=5u
        MP287 N$6180 CK VDD VDD p L=2u W=5u
        MN293 N$6169 N$6173 N$6170 GND n L=2u W=6u
        MN260 N$6201 CK GND GND n L=2u W=5u
        MP260 N$6201 CK VDD VDD p L=2u W=5u
        MN259 N$6196 N$6198 GND GND n L=2u W=6u
        MP412 N$6616 N$6621 VDD VDD p L=2u W=3u
        MP411 N$6619 N$6622 VDD VDD p L=2u W=3u
        MN416 N$6610 N$6624 GND GND n L=2u W=3u
        MN415 N$6611 N$6625 N$6610 GND n L=2u W=3u
        MN263 N$6192 N$6195 GND GND n L=2u W=6u
        MP263 N$6192 N$6195 VDD VDD p L=2u W=6u
        MP262 N$6195 N$6194 N$6193 VDD p L=2u W=6u
        MN262 N$6193 CK N$6195 GND n L=2u W=6u
        MP417 N$6613 N$6621 N$6614 VDD p L=2u W=3u
        MP416 N$6614 N$6624 N$6615 VDD p L=2u W=3u
        MP420 N$6606 N$6605 VDD VDD p L=2u W=3u
        MP266 N$6191 CK N$6190 VDD p L=2u W=6u
        MN298 N$6165 CK N$6167 GND n L=2u W=6u
        MP297 N$5065 CK N$6167 VDD p L=2u W=6u
        MN265 N$6191 CK N$6193 GND n L=2u W=6u
        MP302 N$6163 CK N$6162 VDD p L=2u W=6u
        MN302 N$6162 N$6166 N$6163 GND n L=2u W=6u
        MP301 N$6165 N$6166 N$6163 VDD p L=2u W=6u
        MN301 N$6163 CK N$6165 GND n L=2u W=6u
        MN300 N$6165 N$6164 GND GND n L=2u W=6u
        MP300 N$6165 N$6164 VDD VDD p L=2u W=6u
        MN306 N$6160 N$6159 N$5069 GND n L=2u W=6u
        MN305 N$6166 CK GND GND n L=2u W=5u
        MP305 N$6166 CK VDD VDD p L=2u W=5u
        MN304 N$6161 N$6163 GND GND n L=2u W=6u
        MP304 N$6161 N$6163 VDD VDD p L=2u W=6u
        MN303 N$6162 N$6161 GND GND n L=2u W=6u
        MP303 N$6162 N$6161 VDD VDD p L=2u W=6u
        MP309 N$6158 N$6157 VDD VDD p L=2u W=6u
        MP276 N$6183 N$6182 VDD VDD p L=2u W=6u
        MP275 N$6184 CK N$6183 VDD p L=2u W=6u
        MN275 N$6183 N$6187 N$6184 GND n L=2u W=6u
        MN166 N$6209 N$6208 N$5073 GND n L=2u W=6u
        MN165 N$6217 CK GND GND n L=2u W=5u
        MP248 N$6205 CK N$6204 VDD p L=2u W=6u
        MN248 N$6204 N$6208 N$6205 GND n L=2u W=6u
        MP279 N$5057 CK N$6181 VDD p L=2u W=6u
        MN279 N$6181 N$6180 N$5057 GND n L=2u W=6u
        MN278 N$6187 CK GND GND n L=2u W=5u
        MP278 N$6187 CK VDD VDD p L=2u W=5u
        MN168 N$6206 N$6209 GND GND n L=2u W=6u
        MN251 N$6208 CK GND GND n L=2u W=5u
        MP251 N$6208 CK VDD VDD p L=2u W=5u
        MN282 N$6179 N$6178 GND GND n L=2u W=6u
        MP331 GND N$6151 N$6930 VDD p L=2u W=5u
        MN330 N$6931 N$6151 N$6169 GND n L=2u W=5u
        MP281 N$6178 N$6181 VDD VDD p L=2u W=6u
        MP313 N$6154 N$6156 VDD VDD p L=2u W=6u
        MP318 GND N$6151 N$6921 VDD p L=2u W=5u
        MN317 N$6151 N$8380 GND GND n L=2u W=5u
        MP317 N$6151 N$8380 VDD VDD p L=2u W=5u
        MN316 N$6221 N$6151 N$6211 GND n L=2u W=5u
        MP316 N$6211 N$8380 N$6221 VDD p L=2u W=5u
        MN315 N$6221 N$8380 GND GND n L=2u W=5u
        MP315 GND N$6151 N$6221 VDD p L=2u W=5u
        MP321 N$6197 N$8380 N$6922 VDD p L=2u W=5u
        MN320 N$6922 N$8380 GND GND n L=2u W=5u
        MP320 GND N$6151 N$6922 VDD p L=2u W=5u
        MN319 N$6921 N$6151 N$6204 GND n L=2u W=5u
        MP319 N$6204 N$8380 N$6921 VDD p L=2u W=5u
        MP292 N$6172 N$6173 N$6170 VDD p L=2u W=6u
        MN292 N$6170 CK N$6172 GND n L=2u W=6u
        MN291 N$6172 N$6171 GND GND n L=2u W=6u
        MP259 N$6196 N$6198 VDD VDD p L=2u W=6u
        MN258 N$6197 N$6196 GND GND n L=2u W=6u
        MN264 N$6193 N$6192 GND GND n L=2u W=6u
        MP264 N$6193 N$6192 VDD VDD p L=2u W=6u
        MN295 N$6168 N$6170 GND GND n L=2u W=6u
        MP295 N$6168 N$6170 VDD VDD p L=2u W=6u
        MN294 N$6169 N$6168 GND GND n L=2u W=6u
        MP294 N$6169 N$6168 VDD VDD p L=2u W=6u
        MP261 N$5049 CK N$6195 VDD p L=2u W=6u
        MN267 N$6190 N$6189 GND GND n L=2u W=6u
        MP267 N$6190 N$6189 VDD VDD p L=2u W=6u
        MP298 N$6167 N$6166 N$6165 VDD p L=2u W=6u
        MP134 N$3358 N$6933 N$5049 VDD p L=2u W=5u
        MN313 N$6154 N$6156 GND GND n L=2u W=6u
        MN339 N$6250 N$6933 N$6922 GND n L=2u W=5u
        MP339 N$6922 N$8380 N$6250 VDD p L=2u W=5u
        MN338 N$6248 N$8380 N$6204 GND n L=2u W=5u
        MN347 N$6259 N$6933 N$6931 GND n L=2u W=5u
        MP347 N$6931 N$8380 N$6259 VDD p L=2u W=5u
        MN346 N$6257 N$8380 N$6176 GND n L=2u W=5u
        MP346 N$6176 N$6933 N$6257 VDD p L=2u W=5u
        MN345 N$6257 N$6933 N$6925 GND n L=2u W=5u
        MP345 N$6925 N$8380 N$6257 VDD p L=2u W=5u
        MN350 N$6261 N$8380 N$6162 GND n L=2u W=5u
        MP350 N$6162 N$6933 N$6261 VDD p L=2u W=5u
        MN349 N$6261 N$6933 N$6930 GND n L=2u W=5u
        MP349 N$6930 N$8380 N$6261 VDD p L=2u W=5u
        MN348 N$6259 N$8380 N$6169 GND n L=2u W=5u
        MN318 N$6921 N$8380 GND GND n L=2u W=5u
        MN324 N$6924 N$8380 GND GND n L=2u W=5u
        MP324 GND N$6151 N$6924 VDD p L=2u W=5u
        MP274 N$6186 N$6187 N$6184 VDD p L=2u W=6u
        MN274 N$6184 CK N$6186 GND n L=2u W=6u
        MP280 N$6181 N$6180 N$6179 VDD p L=2u W=6u
        MN280 N$6179 CK N$6181 GND n L=2u W=6u
        MN321 N$6922 N$6151 N$6197 GND n L=2u W=5u
        MN328 N$6925 N$6151 N$6176 GND n L=2u W=5u
        MP328 N$6176 N$8380 N$6925 VDD p L=2u W=5u
        MN327 N$6925 N$8380 GND GND n L=2u W=5u
        MN277 N$6182 N$6184 GND GND n L=2u W=6u
        MP283 N$6179 N$6180 N$6177 VDD p L=2u W=6u
        MN283 N$6177 CK N$6179 GND n L=2u W=6u
        MN331 N$6930 N$8380 GND GND n L=2u W=5u
        MP141 N$6678 N$6683 VDD VDD p L=2u W=6u
        MN141 N$6678 N$6683 GND GND n L=2u W=6u
        MN135 N$6681 N$6678 GND GND n L=2u W=6u
        MN132 N$6676 N$9207 N$6681 GND n L=2u W=6u
        MN129 N$6680 N$6683 GND GND n L=2u W=6u
        MN126 N$6676 N$6677 N$6680 GND n L=2u W=6u
        MP135 N$6676 N$6683 N$6675 VDD p L=2u W=6u
        MP132 N$6675 N$6678 VDD VDD p L=2u W=6u
        MP129 N$6676 N$6677 N$6675 VDD p L=2u W=6u
        MN125 N$5486 N$6668 GND GND n L=2u W=5u
        MP125 N$5486 N$6668 VDD VDD p L=2u W=5u
        MN124 N$6668 N$6664 GND GND n L=2u W=5u
        MN123 N$6668 N$6662 GND GND n L=2u W=5u
        MN122 N$6668 N$6660 GND GND n L=2u W=5u
        MN121 N$6668 N$6659 GND GND n L=2u W=5u
        MP124 N$6668 N$6664 N$6667 VDD p L=2u W=5u
        MP123 N$6667 N$6662 N$6666 VDD p L=2u W=5u
        MP122 N$6666 N$6660 N$6665 VDD p L=2u W=5u
        MN323 N$6923 N$6151 N$6190 GND n L=2u W=5u
        MP323 N$6190 N$8380 N$6923 VDD p L=2u W=5u
        MN322 N$6923 N$8380 GND GND n L=2u W=5u
        MP322 GND N$6151 N$6923 VDD p L=2u W=5u
        MP121 N$6665 N$6659 VDD VDD p L=2u W=5u
        MP327 GND N$6151 N$6925 VDD p L=2u W=5u
        MN325 N$6924 N$6151 N$6183 GND n L=2u W=5u
        MP325 N$6183 N$8380 N$6924 VDD p L=2u W=5u
        MP151 N$6102 N$6651 N$5078 VDD p L=2u W=5u
        MP354 N$6246 N$6689 N$6235 VDD p L=2u W=5u
        MN56 N$1726 N$1722 GND GND n L=2u W=3u
        MN52 N$1724 N$6243 N$1725 GND n L=2u W=3u
        MP130 N$1709 N$6651 N$5045 VDD p L=2u W=5u
        MN130 N$5045 N$6933 N$1709 GND n L=2u W=5u
        MP29 N$1693 N$6233 VDD VDD p L=2u W=3u
        MN144 N$6682 N$6676 GND GND n L=2u W=6u
        MP144 N$6682 N$6676 VDD VDD p L=2u W=6u
        MN138 N$6677 N$9207 GND GND n L=2u W=6u
        MP138 N$6677 N$9207 VDD VDD p L=2u W=6u
        MP694 N$6358 N$6359 N$6356 VDD p L=2u W=6u
        MP700 N$6354 N$6353 N$6352 VDD p L=2u W=6u
        MN667 N$6470 N$6376 N$6485 GND n L=2u W=5u
        MP667 N$6485 N$6515 N$6470 VDD p L=2u W=5u
        MN666 N$6470 N$6515 N$6444 GND n L=2u W=5u
        MP672 N$9216 N$6376 N$9221 VDD p L=2u W=5u
        MP698 N$6359 CK VDD VDD p L=2u W=5u
        MN697 N$6355 N$6356 GND GND n L=2u W=6u
        MP703 N$6352 N$6353 N$6350 VDD p L=2u W=6u
        MN670 N$6454 N$6515 N$6442 GND n L=2u W=5u
        MP670 N$6442 N$6376 N$6454 VDD p L=2u W=5u
        MN669 N$6462 N$6376 N$6484 GND n L=2u W=5u
        MN701 N$6351 N$6354 GND GND n L=2u W=6u
        MN695 N$6269 N$6359 N$6356 GND n L=2u W=6u
        MP695 N$6356 CK N$6269 VDD p L=2u W=6u
        MN673 N$9221 N$6376 GND GND n L=2u W=5u
        MP673 GND N$6515 N$9221 VDD p L=2u W=5u
        MN672 N$9221 N$6515 N$9216 GND n L=2u W=5u
        MN678 N$6369 N$6376 GND GND n L=2u W=5u
        MP678 GND N$6515 N$6369 VDD p L=2u W=5u
        MN677 N$6369 N$6515 N$6393 GND n L=2u W=5u
        MP677 N$6393 N$6376 N$6369 VDD p L=2u W=5u
        MN676 N$6370 N$6376 GND GND n L=2u W=5u
        MP676 GND N$6515 N$6370 VDD p L=2u W=5u
        MN675 N$6370 N$6515 N$6408 GND n L=2u W=5u
        MP681 N$9221 CK N$6366 VDD p L=2u W=6u
        MN681 N$6366 N$9223 N$9221 GND n L=2u W=6u
        MN680 N$6368 N$6376 GND GND n L=2u W=5u
        MP662 N$6406 N$6443 VDD VDD p L=2u W=3u
        MN661 N$6391 N$6442 GND GND n L=2u W=3u
        MP661 N$6391 N$6442 VDD VDD p L=2u W=3u
        MN660 N$6421 N$6444 GND GND n L=2u W=3u
        MP666 N$6444 N$6376 N$6470 VDD p L=2u W=5u
        MN665 N$6376 N$6515 GND GND n L=2u W=5u
        MP665 N$6376 N$6515 VDD VDD p L=2u W=5u
        MN664 N$6479 N$6376 N$6487 GND n L=2u W=5u
        MP664 N$6487 N$6515 N$6479 VDD p L=2u W=5u
        MN870 N$8378 N$8379 GND GND n L=2u W=5u
        MP870 N$8378 N$8379 VDD VDD p L=2u W=5u
        MN869 N$8379 N$8380 GND GND n L=2u W=5u
        MN868 N$8379 N$6658 GND GND n L=2u W=5u
        MP869 N$8379 N$8380 N$8375 VDD p L=2u W=5u
        MP868 N$8375 N$6658 VDD VDD p L=2u W=5u
        MN867 N$7766 N$8173 N$8378 GND n L=2u W=5u
        MP867 N$8378 N$6499 N$7766 VDD p L=2u W=5u
        MN866 N$7766 N$6499 N$6658 GND n L=2u W=5u
        MP866 N$6658 N$8173 N$7766 VDD p L=2u W=5u
        MP370 N$6947 N$6913 N$6896 VDD p L=2u W=5u
        MN662 N$6406 N$6443 GND GND n L=2u W=3u
        MP663 N$9213 N$6376 N$6479 VDD p L=2u W=5u
        MN657 N$6382 N$6403 N$6380 GND n L=2u W=3u
        MP658 N$6378 N$6382 VDD VDD p L=2u W=3u
        MN599 N$6443 N$6515 N$6490 GND n L=2u W=5u
        MP599 N$6490 N$6447 N$6443 VDD p L=2u W=5u
        MN598 N$6444 N$6447 GND GND n L=2u W=5u
        MP598 GND N$6515 N$6444 VDD p L=2u W=5u
        MN597 N$6444 N$6515 N$6526 GND n L=2u W=5u
        MP597 N$6526 N$6447 N$6444 VDD p L=2u W=5u
        MN620 N$6416 N$6421 GND GND n L=2u W=3u
        MN602 N$6442 N$6447 GND GND n L=2u W=5u
        MP602 GND N$6515 N$6442 VDD p L=2u W=5u
        MN601 N$6442 N$6515 N$6519 GND n L=2u W=5u
        MP601 N$6519 N$6447 N$6442 VDD p L=2u W=5u
        MN600 N$6443 N$6447 GND GND n L=2u W=5u
        MN618 N$6417 H1 GND GND n L=2u W=3u
        MN619 N$6419 N$8383 N$6417 GND n L=2u W=3u
        MP616 N$9216 N$8594 VDD VDD p L=2u W=3u
        MN615 N$8594 C0 N$8596 GND n L=2u W=3u
        MN614 N$8594 N$8588 N$8595 GND n L=2u W=3u
        MN613 N$8597 N$8586 GND GND n L=2u W=3u
        MN612 N$8596 H0 N$8597 GND n L=2u W=3u
        MN611 N$8595 C0 GND GND n L=2u W=3u
        MN610 N$8595 N$8586 GND GND n L=2u W=3u
        MP600 GND N$6515 N$6443 VDD p L=2u W=5u
        MP549 N$6494 N$6488 N$6487 VDD p L=2u W=5u
        MN549 N$6487 N$6499 N$6494 GND n L=2u W=5u
        MP550 GND N$6499 N$6487 VDD p L=2u W=5u
        MP548 N$6490 RST N$6588 VDD p L=2u W=5u
        MN553 N$6485 N$6488 GND GND n L=2u W=5u
        MP553 GND N$6499 N$6485 VDD p L=2u W=5u
        MN578 N$6460 N$6464 GND GND n L=2u W=6u
        MP552 N$6533 N$6488 N$6485 VDD p L=2u W=5u
        MP495 N$6527 CK N$6526 VDD p L=2u W=6u
        MP536 N$9207 N$6658 VDD VDD p L=2u W=6u
        MP500 N$6524 N$6523 N$6522 VDD p L=2u W=6u
        MN500 N$6522 CK N$6524 GND n L=2u W=6u
        MP499 N$6547 CK N$6524 VDD p L=2u W=6u
        MN499 N$6524 N$6523 N$6547 GND n L=2u W=6u
        MN498 N$6530 CK GND GND n L=2u W=5u
        MP498 N$6530 CK VDD VDD p L=2u W=5u
        MN504 N$6519 N$6523 N$6520 GND n L=2u W=6u
        MP503 N$6522 N$6523 N$6520 VDD p L=2u W=6u
        MN503 N$6520 CK N$6522 GND n L=2u W=6u
        MN502 N$6522 N$6521 GND GND n L=2u W=6u
        MP502 N$6522 N$6521 VDD VDD p L=2u W=6u
        MN501 N$6521 N$6524 GND GND n L=2u W=6u
        MP501 N$6521 N$6524 VDD VDD p L=2u W=6u
        MP507 N$6523 CK VDD VDD p L=2u W=5u
        MN506 N$6518 N$6520 GND GND n L=2u W=6u
        MP506 N$6518 N$6520 VDD VDD p L=2u W=6u
        MN505 N$6519 N$6518 GND GND n L=2u W=6u
        MP546 N$6526 RST N$6605 VDD p L=2u W=5u
        MN545 N$6605 RST GND GND n L=2u W=5u
        MP545 GND N$6497 N$6605 VDD p L=2u W=5u
        MN550 N$6487 N$6488 GND GND n L=2u W=5u
        MN517 N$6515 N$6516 GND GND n L=2u W=5u
        MP518 N$6515 N$6658 N$6517 VDD p L=2u W=5u
        MP517 N$6517 N$6516 VDD VDD p L=2u W=5u
        MN507 N$6523 CK GND GND n L=2u W=5u
        MP496 N$6526 N$6525 VDD VDD p L=2u W=6u
        MN548 N$6588 N$6497 N$6490 GND n L=2u W=5u
        MP521 N$6550 CK N$6510 VDD p L=2u W=6u
        MP78 N$1755 N$6255 VDD VDD p L=2u W=3u
        MN197 N$6277 N$6542 GND GND n L=2u W=3u
        MP769 N$6278 N$6284 N$6281 VDD p L=2u W=3u
        MP768 N$6278 C0 N$6279 VDD p L=2u W=3u
        MP201 N$6279 N$6286 N$6280 VDD p L=2u W=3u
        MN770 N$6554 N$6278 GND GND n L=2u W=3u
        MP770 N$6554 N$6278 VDD VDD p L=2u W=3u
        MN769 N$6278 C0 N$6276 GND n L=2u W=3u
        MN768 N$6278 N$6284 N$6277 GND n L=2u W=3u
        MN201 N$6275 N$6286 GND GND n L=2u W=3u
        MN200 N$6276 N$6542 N$6275 GND n L=2u W=3u
        MP773 N$6519 RST N$6572 VDD p L=2u W=5u
        MN772 N$6572 RST GND GND n L=2u W=5u
        MP772 GND N$6497 N$6572 VDD p L=2u W=5u
        MN771 N$6286 H0 GND GND n L=2u W=3u
        MP7 N$231 GND VDD VDD p L=2u W=3u
        MP60 N$1732 N$1489 N$1728 VDD p L=2u W=3u
        MP59 N$1731 N$6225 N$1728 VDD p L=2u W=3u
        MN87 N$1768 N$1752 N$1771 GND n L=2u W=3u
        MN199 N$6277 C0 GND GND n L=2u W=3u
        MN195 N$6283 N$6286 GND GND n L=2u W=3u
        MN15 N$1276 N$1274 GND GND n L=2u W=3u
        MP111 N$1794 N$1786 N$1791 VDD p L=2u W=3u
        MP110 N$1794 N$1770 N$1793 VDD p L=2u W=3u
        MP109 N$1793 N$4416 N$1792 VDD p L=2u W=3u
        MP31 N$1696 GND N$1693 VDD p L=2u W=3u
        MN449 N$6567 N$6572 GND GND n L=2u W=3u
        MN485 N$6534 CK N$6536 GND n L=2u W=6u
        MP452 N$6569 N$6572 N$6570 VDD p L=2u W=3u
        MP451 N$6569 N$6584 N$6573 VDD p L=2u W=3u
        MP450 N$6570 N$6571 N$6573 VDD p L=2u W=3u
        MP455 N$6565 N$6572 VDD VDD p L=2u W=3u
        MP454 N$6565 N$6584 VDD VDD p L=2u W=3u
        MP453 N$6683 N$6569 VDD VDD p L=2u W=3u
        MN453 N$6569 N$6572 N$6566 GND n L=2u W=3u
        MN452 N$6567 N$6571 GND GND n L=2u W=3u
        MN451 N$6566 N$6571 GND GND n L=2u W=3u
        MN455 N$6561 N$6571 GND GND n L=2u W=3u
        MN454 N$6561 N$6572 GND GND n L=2u W=3u
        MP460 N$6562 N$6569 N$6565 VDD p L=2u W=3u
        MP459 N$6562 N$6584 N$6563 VDD p L=2u W=3u
        MP458 N$6563 N$6571 N$6564 VDD p L=2u W=3u
        MP457 N$6564 N$6572 N$6565 VDD p L=2u W=3u
        MP456 N$6565 N$6571 VDD VDD p L=2u W=3u
        MP489 N$6539 CK VDD VDD p L=2u W=5u
        MN488 N$6532 N$6534 GND GND n L=2u W=6u
        MP494 N$6529 N$6530 N$6527 VDD p L=2u W=6u
        MN494 N$6527 CK N$6529 GND n L=2u W=6u
        MN457 N$6560 N$6572 N$6559 GND n L=2u W=3u
        MN456 N$6561 N$6584 GND GND n L=2u W=3u
        MP464 N$6571 GND VDD VDD p L=2u W=3u
        MN463 N$6604 H2 GND GND n L=2u W=3u
        MN497 N$6525 N$6527 GND GND n L=2u W=6u
        MP497 N$6525 N$6527 VDD VDD p L=2u W=6u
        MN450 N$6569 N$6584 N$6567 GND n L=2u W=3u
        MN568 N$6469 CK N$6472 GND n L=2u W=6u
        MN575 N$6471 CK GND GND n L=2u W=5u
        MP581 N$6459 CK N$6911 VDD p L=2u W=6u
        MN581 N$6911 N$6463 N$6459 GND n L=2u W=6u
        MP580 N$6461 N$6463 N$6459 VDD p L=2u W=6u
        MN580 N$6459 CK N$6461 GND n L=2u W=6u
        MN579 N$6461 N$6460 GND GND n L=2u W=6u
        MP579 N$6461 N$6460 VDD VDD p L=2u W=6u
        MN576 N$6464 N$6463 N$6462 GND n L=2u W=6u
        MN207 N$6919 N$6904 GND GND n L=2u W=5u
        MP584 N$6463 CK VDD VDD p L=2u W=5u
        MN583 N$6457 N$6459 GND GND n L=2u W=6u
        MP583 N$6457 N$6459 VDD VDD p L=2u W=6u
        MN582 N$6911 N$6457 GND GND n L=2u W=6u
        MP582 N$6911 N$6457 VDD VDD p L=2u W=6u
        MP615 N$8594 N$8588 N$8591 VDD p L=2u W=3u
        MP614 N$8594 C0 N$8593 VDD p L=2u W=3u
        MP613 N$8593 N$8586 N$8592 VDD p L=2u W=3u
        MP612 N$8592 H0 N$8591 VDD p L=2u W=3u
        MP611 N$8591 N$8586 VDD VDD p L=2u W=3u
        MP610 N$8591 H0 VDD VDD p L=2u W=3u
        MP609 N$8591 C0 VDD VDD p L=2u W=3u
        MP608 N$8383 N$8588 VDD VDD p L=2u W=3u
        MN608 N$8588 H0 N$8590 GND n L=2u W=3u
        MN607 N$8589 N$8586 GND GND n L=2u W=3u
        MN606 N$8590 N$8586 GND GND n L=2u W=3u
        MN605 N$8588 C0 N$8589 GND n L=2u W=3u
        MN604 N$8589 H0 GND GND n L=2u W=3u
        MN603 N$8383 N$8588 GND GND n L=2u W=3u
        MP607 N$8588 H0 N$8587 VDD p L=2u W=3u
        MP606 N$8588 C0 N$8585 VDD p L=2u W=3u
        MN214 N$6916 N$7766 GND GND n L=2u W=5u
        MP214 GND N$6904 N$6916 VDD p L=2u W=5u
        MN213 N$6916 N$6904 A1 GND n L=2u W=5u
        MP213 A1 N$7766 N$6916 VDD p L=2u W=5u
        MN224 N$6914 N$6905 N$6919 GND n L=2u W=5u
        MP212 GND N$6904 N$6917 VDD p L=2u W=5u
        MN211 N$6917 N$6904 A2 GND n L=2u W=5u
        MP211 A2 N$7766 N$6917 VDD p L=2u W=5u
        MN210 N$6918 N$7766 GND GND n L=2u W=5u
        MP210 GND N$6904 N$6918 VDD p L=2u W=5u
        MN209 N$6918 N$6904 A3 GND n L=2u W=5u
        MP209 A3 N$7766 N$6918 VDD p L=2u W=5u
        MN212 N$6917 N$7766 GND GND n L=2u W=5u
        MP215 A0 N$7766 N$6915 VDD p L=2u W=5u
        MN208 N$6919 N$7766 GND GND n L=2u W=5u
        MP208 GND N$6904 N$6919 VDD p L=2u W=5u
        MP403 N$6769 N$6696 N$6768 VDD p L=2u W=3u
        MP402 N$6768 N$6921 N$6767 VDD p L=2u W=3u
        MP401 N$6767 N$6696 VDD VDD p L=2u W=3u
        MP371 N$6948 N$6911 N$6883 VDD p L=2u W=5u
        MP380 N$6745 N$6900 VDD VDD p L=2u W=3u
        MN370 N$6896 N$6911 N$6947 GND n L=2u W=5u
        MP404 N$6770 N$6749 N$6769 VDD p L=2u W=3u
        MN397 N$6765 N$6696 GND GND n L=2u W=3u
        MN396 N$6766 N$6696 GND GND n L=2u W=3u
        MN395 N$6762 N$6749 N$6765 GND n L=2u W=3u
        MN351 N$6895 N$6911 N$6948 GND n L=2u W=5u
        MP329 GND N$6151 N$6931 VDD p L=2u W=5u
        MN333 OUT8 N$6151 N$6633 GND n L=2u W=5u
        MN326 OUT8 N$8380 GND GND n L=2u W=5u
        MP326 GND N$6151 OUT8 VDD p L=2u W=5u
        MN332 N$6930 N$6151 N$6162 GND n L=2u W=5u
        MP332 N$6162 N$8380 N$6930 VDD p L=2u W=5u
        MP335 N$6211 N$6933 N$6246 VDD p L=2u W=5u
        MN334 N$6246 N$6933 N$6221 GND n L=2u W=5u
        MP334 N$6221 N$8380 N$6246 VDD p L=2u W=5u
        MN329 N$6931 N$8380 GND GND n L=2u W=5u
        MN297 N$6167 N$6166 N$5065 GND n L=2u W=6u
        MN308 N$6157 N$6160 GND GND n L=2u W=6u
        MP308 N$6157 N$6160 VDD VDD p L=2u W=6u
        MP307 N$6160 N$6159 N$6158 VDD p L=2u W=6u
        MN307 N$6158 CK N$6160 GND n L=2u W=6u
        MP306 N$5069 CK N$6160 VDD p L=2u W=6u
        MN312 N$6633 N$6154 GND GND n L=2u W=6u
        MN352 N$6896 N$6913 N$6914 GND n L=2u W=5u
        MP851 N$6884 S3 VDD VDD p L=2u W=5u
        MN865 N$6900 S3 GND GND n L=2u W=5u
        MN850 N$6891 S3 N$6896 GND n L=2u W=5u
        MN218 N$6730 N$6910 N$6864 GND n L=2u W=5u
        MP218 N$6864 N$6905 N$6730 VDD p L=2u W=5u
        MN217 N$6730 N$6905 N$6714 GND n L=2u W=5u
        MP379 N$6745 N$6221 VDD VDD p L=2u W=3u
        MP203 GND N$7766 N$6864 VDD p L=2u W=5u
        MN202 N$6904 N$7766 GND GND n L=2u W=5u
        MP202 N$6904 N$7766 VDD VDD p L=2u W=5u
        MP333 N$6633 N$8380 OUT8 VDD p L=2u W=5u
        MN851 N$6884 S3 GND GND n L=2u W=5u
        MN150 N$6714 N$7766 GND GND n L=2u W=5u
        MP150 GND N$6904 N$6714 VDD p L=2u W=5u
        MN147 N$6714 N$6904 GND GND n L=2u W=5u
        MN100 N$1789 N$6244 GND GND n L=2u W=3u
        MP36 N$1702 N$6233 VDD VDD p L=2u W=3u
        MP72 N$1746 N$6223 VDD VDD p L=2u W=3u
        MP99 N$1782 N$6244 VDD VDD p L=2u W=3u
        MP100 N$1782 N$4416 VDD VDD p L=2u W=3u
        MP92 N$1773 N$6238 VDD VDD p L=2u W=3u
        MN101 N$1786 N$1770 N$1789 GND n L=2u W=3u
        MP139 N$1762 N$6651 N$5057 VDD p L=2u W=5u
        MN37 N$1706 N$1276 GND GND n L=2u W=3u
        MN143 N$5061 N$6651 N$1798 GND n L=2u W=5u
        MP143 N$1798 N$6933 N$5061 VDD p L=2u W=5u
        MN137 N$5053 N$6651 N$1762 GND n L=2u W=5u
        MP137 N$1762 N$6933 N$5053 VDD p L=2u W=5u
        MN136 N$5053 N$6933 N$3358 GND n L=2u W=5u
        MP136 N$3358 N$6651 N$5053 VDD p L=2u W=5u
        MP68 N$1740 N$1489 N$1739 VDD p L=2u W=3u
        MN75 N$1753 N$6223 GND GND n L=2u W=3u
        MN153 N$6651 N$6933 GND GND n L=2u W=5u
        MP153 N$6651 N$6933 VDD VDD p L=2u W=5u
        MN151 N$5078 N$6933 N$6102 GND n L=2u W=5u
        MN39 N$1708 GND GND GND n L=2u W=3u
        MP149 GND N$6933 N$5069 VDD p L=2u W=5u
        MP85 N$1764 N$6238 VDD VDD p L=2u W=3u
        MP140 N$1780 N$6933 N$5057 VDD p L=2u W=5u
        MN35 N$1706 N$6233 GND GND n L=2u W=3u
        MN72 N$1753 N$6255 GND GND n L=2u W=3u
        MN154 N$6232 N$5486 GND GND n L=2u W=5u
        MP155 N$6232 GND N$5485 VDD p L=2u W=5u
        MP154 N$5485 N$5486 VDD VDD p L=2u W=5u
        MN357 N$6234 N$6266 N$6248 GND n L=2u W=5u
        MN164 N$6210 N$6212 GND GND n L=2u W=6u
        MP164 N$6210 N$6212 VDD VDD p L=2u W=6u
        MN163 N$6211 N$6210 GND GND n L=2u W=6u
        MP163 N$6211 N$6210 VDD VDD p L=2u W=6u
        MP162 N$6212 CK N$6211 VDD p L=2u W=6u
        MN162 N$6211 N$6217 N$6212 GND n L=2u W=6u
        MP168 N$6206 N$6209 VDD VDD p L=2u W=6u
        MP56 N$1726 N$1722 VDD VDD p L=2u W=3u
        MP159 N$6213 N$6218 VDD VDD p L=2u W=6u
        MN159 N$6213 N$6218 GND GND n L=2u W=6u
        MP344 N$6183 N$6933 N$6254 VDD p L=2u W=5u
        MN343 N$6254 N$6933 N$6924 GND n L=2u W=5u
        MP343 N$6924 N$8380 N$6254 VDD p L=2u W=5u
        MN342 N$6252 N$8380 N$6190 GND n L=2u W=5u
        MN344 N$6254 N$8380 N$6183 GND n L=2u W=5u
        MP342 N$6190 N$6933 N$6252 VDD p L=2u W=5u
        MP245 GND N$5896 N$4416 VDD p L=2u W=6u
        MP362 GND N$6266 N$6236 VDD p L=2u W=5u
        MN363 N$6236 N$6266 N$6254 GND n L=2u W=5u
        MN361 N$6243 N$6266 N$6252 GND n L=2u W=5u
        MP361 N$6252 N$6689 N$6243 VDD p L=2u W=5u
        MN90 N$1768 N$6238 N$1772 GND n L=2u W=3u
        MN369 N$6244 N$6266 N$6261 GND n L=2u W=5u
        MP369 N$6261 N$6689 N$6244 VDD p L=2u W=5u
        MN368 N$6244 N$6689 GND GND n L=2u W=5u
        MP363 N$6254 N$6689 N$6236 VDD p L=2u W=5u
        MN7 N$239 N$6235 GND GND n L=2u W=3u
        MP98 N$1780 N$1776 VDD VDD p L=2u W=3u
        MN366 N$6238 N$6689 GND GND n L=2u W=5u
        MP147 GND N$7766 N$6714 VDD p L=2u W=5u
        MN86 N$1771 N$6238 GND GND n L=2u W=3u
        MN85 N$1770 N$1768 GND GND n L=2u W=3u
        MP89 N$1768 N$6238 N$1767 VDD p L=2u W=3u
        MP88 N$1768 N$1752 N$1764 VDD p L=2u W=3u
        MP87 N$1767 N$4413 N$1764 VDD p L=2u W=3u
        MP86 N$1764 N$4413 VDD VDD p L=2u W=3u
        MN84 N$1762 N$1758 GND GND n L=2u W=3u
        MP84 N$1762 N$1758 VDD VDD p L=2u W=3u
        MN83 N$1758 N$1734 N$1760 GND n L=2u W=3u
        MN82 N$1758 N$1750 N$1759 GND n L=2u W=3u
        MN107 N$1795 N$1770 GND GND n L=2u W=3u
        MN106 N$1795 N$4416 GND GND n L=2u W=3u
        MP243 GND N$5896 N$6223 VDD p L=2u W=6u
        MP37 N$1702 GND VDD VDD p L=2u W=3u
        MN92 N$1777 N$4413 GND GND n L=2u W=3u
        MN152 N$5078 N$6651 N$1286 GND n L=2u W=5u
        MP152 N$1286 N$6933 N$5078 VDD p L=2u W=5u
        MN516 N$6785 N$6764 GND GND n L=2u W=3u
        MN515 N$6785 N$6887 GND GND n L=2u W=3u
        MN514 N$6785 N$6922 GND GND n L=2u W=3u
        MP777 N$6784 N$6777 N$6781 VDD p L=2u W=3u
        MP47 N$1715 N$6243 N$1714 VDD p L=2u W=3u
        MP63 N$1737 N$1489 VDD VDD p L=2u W=3u
        MN155 N$6232 GND GND GND n L=2u W=5u
        MP515 N$6781 N$6922 VDD VDD p L=2u W=3u
        MP514 N$6781 N$6764 VDD VDD p L=2u W=3u
        MP513 N$6865 N$6777 VDD VDD p L=2u W=3u
        MN47 N$1717 GND GND GND n L=2u W=3u
        MN858 N$6888 N$6884 N$6883 GND n L=2u W=5u
        MP858 N$6883 S3 N$6888 VDD p L=2u W=5u
        MN857 N$6889 S3 N$6956 GND n L=2u W=5u
        MP857 N$6956 N$6884 N$6889 VDD p L=2u W=5u
        MN856 N$6889 N$6884 N$6896 GND n L=2u W=5u
        MP856 N$6896 S3 N$6889 VDD p L=2u W=5u
        MN855 N$6867 S3 N$6957 GND n L=2u W=5u
        MP855 N$6957 N$6884 N$6867 VDD p L=2u W=5u
        MN854 N$6867 N$6884 N$6895 GND n L=2u W=5u
        MP854 N$6895 S3 N$6867 VDD p L=2u W=5u
        MN853 N$6890 S3 N$6883 GND n L=2u W=5u
        MP853 N$6883 N$6884 N$6890 VDD p L=2u W=5u
        MN852 N$6890 N$6884 N$6894 GND n L=2u W=5u
        MP852 N$6894 S3 N$6890 VDD p L=2u W=5u
        MP205 GND N$7766 N$6920 VDD p L=2u W=5u
        MP311 N$6156 CK N$6633 VDD p L=2u W=6u
        MN311 N$6633 N$6159 N$6156 GND n L=2u W=6u
        MP310 N$6158 N$6159 N$6156 VDD p L=2u W=6u
        MN205 N$6920 N$6904 GND GND n L=2u W=5u
        MP312 N$6633 N$6154 VDD VDD p L=2u W=6u
        MP860 N$6957 S3 N$6887 VDD p L=2u W=5u
        MN859 N$6888 S3 N$6955 GND n L=2u W=5u
        MP859 N$6955 N$6884 N$6888 VDD p L=2u W=5u
        MP314 N$6159 CK VDD VDD p L=2u W=5u
        MN228 N$6947 N$6905 N$6917 GND n L=2u W=5u
        MP228 N$6917 N$6910 N$6947 VDD p L=2u W=5u
        MN227 N$6948 N$6910 N$6917 GND n L=2u W=5u
        MP227 N$6917 N$6905 N$6948 VDD p L=2u W=5u
        MP356 GND N$6266 N$6234 VDD p L=2u W=5u
        MN353 N$6235 N$6689 GND GND n L=2u W=5u
        MP22 N$1279 N$6234 VDD VDD p L=2u W=3u
        MP5 N$245 N$6235 N$212 VDD p L=2u W=3u
        MP4 N$245 GND N$209 VDD p L=2u W=3u
        MP3 N$212 GND N$209 VDD p L=2u W=3u
        MN42 N$1709 N$1705 GND GND n L=2u W=3u
        MP80 N$1756 N$6255 N$1755 VDD p L=2u W=3u
        MP81 N$1757 N$6223 N$1756 VDD p L=2u W=3u
        MP82 N$1758 N$1734 N$1757 VDD p L=2u W=3u
        MN6 N$245 N$6235 N$222 GND n L=2u W=3u
        MN9 N$239 GND GND GND n L=2u W=3u
        MN10 N$241 N$6235 N$236 GND n L=2u W=3u
        MN362 N$6236 N$6689 GND GND n L=2u W=5u
        MN60 N$1736 N$6225 GND GND n L=2u W=3u
        MN156 N$5896 N$6232 GND GND n L=2u W=5u
        MP156 N$5896 N$6232 VDD VDD p L=2u W=5u
        MP242 N$6269 N$6232 N$6223 VDD p L=2u W=6u
        MN242 N$6223 N$5896 N$6269 GND n L=2u W=6u
        MP247 GND N$5896 N$4413 VDD p L=2u W=6u
        MP40 N$1705 N$1276 N$1704 VDD p L=2u W=3u
        MN142 N$5061 N$6933 N$1780 GND n L=2u W=5u
        MP142 N$1780 N$6651 N$5061 VDD p L=2u W=5u
        MN127 N$5073 N$6933 N$1286 GND n L=2u W=5u
        MN29 N$1699 N$1697 GND GND n L=2u W=3u
        MN26 N$1282 N$1274 N$1283 GND n L=2u W=3u
        MP27 N$1282 N$1274 N$1279 VDD p L=2u W=3u
        MN21 N$1283 N$6234 GND GND n L=2u W=3u
        MN140 N$5057 N$6651 N$1780 GND n L=2u W=5u
        MN119 N$6664 N$6691 A3 GND n L=2u W=5u
        MP340 N$6197 N$6933 N$6250 VDD p L=2u W=5u
        MP126 N$6675 N$9207 VDD VDD p L=2u W=6u
        MN148 N$5069 N$6933 N$6634 GND n L=2u W=5u
        MN149 N$5069 N$6651 GND GND n L=2u W=5u
        MP148 N$6634 N$6651 N$5069 VDD p L=2u W=5u
        MN51 N$1723 N$1699 GND GND n L=2u W=3u
        MP67 N$1739 N$6225 N$1738 VDD p L=2u W=3u
        MP66 N$1738 N$6236 N$1737 VDD p L=2u W=3u
        MN120 GND N$6319 N$6664 GND n L=2u W=5u
        MN28 N$1286 N$1282 GND GND n L=2u W=3u
        MP28 N$1286 N$1282 VDD VDD p L=2u W=3u
        MN128 N$5073 N$6651 N$1709 GND n L=2u W=5u
        MN40 N$1705 N$1697 N$1706 GND n L=2u W=3u
        MP30 N$1693 GND VDD VDD p L=2u W=3u
        MN62 N$1732 N$6236 N$1736 GND n L=2u W=3u
        MP291 N$6172 N$6171 VDD VDD p L=2u W=6u
        MN290 N$6171 N$6174 GND GND n L=2u W=6u
        MN296 N$6173 CK GND GND n L=2u W=5u
        MP296 N$6173 CK VDD VDD p L=2u W=5u
        MN27 N$1282 N$5 N$1284 GND n L=2u W=3u
        MP58 N$1728 N$6225 VDD VDD p L=2u W=3u
        MN54 N$1722 N$1715 N$1723 GND n L=2u W=3u
        MN53 N$1725 GND GND GND n L=2u W=3u
        MP293 N$6170 CK N$6169 VDD p L=2u W=6u
        MN299 N$6164 N$6167 GND GND n L=2u W=6u
        MP299 N$6164 N$6167 VDD VDD p L=2u W=6u
        MP131 N$1726 N$6933 N$5045 VDD p L=2u W=5u
        MP1 N$209 N$6235 VDD VDD p L=2u W=3u
        MN364 N$6255 N$6689 GND GND n L=2u W=5u
        MP364 GND N$6266 N$6255 VDD p L=2u W=5u
        MN410 N$6618 N$6624 GND GND n L=2u W=3u
        MN409 N$6617 N$6624 GND GND n L=2u W=3u
        MN408 N$6622 N$6621 N$6618 GND n L=2u W=3u
        MN407 N$6618 N$6625 GND GND n L=2u W=3u
        MP348 N$6169 N$6933 N$6259 VDD p L=2u W=5u
        MN411 N$6622 N$6625 N$6617 GND n L=2u W=3u
        MN70 N$3358 N$1740 GND GND n L=2u W=3u
        MP14 N$6102 N$855 VDD VDD p L=2u W=3u
        MP61 N$1732 N$6236 N$1731 VDD p L=2u W=3u
        MP146 N$6634 N$6933 N$5065 VDD p L=2u W=5u
        MN145 N$5065 N$6933 N$1798 GND n L=2u W=5u
        MP145 N$1798 N$6651 N$5065 VDD p L=2u W=5u
        MN2 N$218 N$6235 GND GND n L=2u W=3u
        MN14 N$6102 N$855 GND GND n L=2u W=3u
        MN3 N$245 GND N$218 GND n L=2u W=3u
        MN365 N$6255 N$6266 N$6257 GND n L=2u W=5u
        MP104 N$6634 N$1786 VDD VDD p L=2u W=3u
        MP128 N$1709 N$6933 N$5073 VDD p L=2u W=5u
        MP101 N$1785 N$4416 N$1782 VDD p L=2u W=3u
        MN236 N$6225 N$6232 GND GND n L=2u W=6u
        MP235 N$6268 N$6232 N$6225 VDD p L=2u W=6u
        MN235 N$6225 N$5896 N$6268 GND n L=2u W=6u
        MP127 N$1286 N$6651 N$5073 VDD p L=2u W=5u
        MN61 N$1735 N$6225 GND GND n L=2u W=3u
        MP366 GND N$6266 N$6238 VDD p L=2u W=5u
        MN247 N$4413 N$6232 GND GND n L=2u W=6u
        MP365 N$6257 N$6689 N$6255 VDD p L=2u W=5u
        MP73 N$1749 N$6223 N$1746 VDD p L=2u W=3u
        MP65 N$1737 N$6225 VDD VDD p L=2u W=3u
        MP8 N$231 N$6235 VDD VDD p L=2u W=3u
        MP9 N$231 GND VDD VDD p L=2u W=3u
        MP10 N$226 N$6235 N$231 VDD p L=2u W=3u
        MP11 N$228 GND N$226 VDD p L=2u W=3u
        MP12 N$855 GND N$228 VDD p L=2u W=3u
        MP91 N$1773 N$1752 VDD VDD p L=2u W=3u
        MP74 N$1750 N$1734 N$1746 VDD p L=2u W=3u
        MN4 N$222 GND GND GND n L=2u W=3u
        MN19 N$1277 GND GND GND n L=2u W=3u
        MN64 N$1741 N$6225 GND GND n L=2u W=3u
        MN65 N$1741 N$1489 GND GND n L=2u W=3u
        MN99 N$6634 N$1786 GND GND n L=2u W=3u
        MN63 N$1741 N$6236 GND GND n L=2u W=3u
        MP69 N$1740 N$1732 N$1737 VDD p L=2u W=3u
        MN5 N$218 GND GND GND n L=2u W=3u
        MP103 N$1786 N$6244 N$1785 VDD p L=2u W=3u
        MP102 N$1786 N$1770 N$1782 VDD p L=2u W=3u
        MP45 N$1714 GND N$1711 VDD p L=2u W=3u
        MP44 N$1711 GND VDD VDD p L=2u W=3u
        MP43 N$1711 N$6243 VDD VDD p L=2u W=3u
        MN12 N$855 N$245 N$239 GND n L=2u W=3u
        MP236 GND N$5896 N$6225 VDD p L=2u W=6u
        MN43 N$1489 N$1715 GND GND n L=2u W=3u
        MP160 N$6214 N$6213 VDD VDD p L=2u W=6u
        MN185 N$6490 N$6293 N$6290 GND n L=2u W=6u
        MP35 N$1702 N$1276 VDD VDD p L=2u W=3u
        MN184 N$6290 CK N$6292 GND n L=2u W=6u
        MN183 N$6292 N$6291 GND GND n L=2u W=6u
        MP183 N$6292 N$6291 VDD VDD p L=2u W=6u
        MP189 N$6542 N$6548 N$6299 VDD p L=2u W=5u
        MN188 N$6293 CK GND GND n L=2u W=5u
        MP188 N$6293 CK VDD VDD p L=2u W=5u
        MN187 N$6289 N$6290 GND GND n L=2u W=6u
        MP187 N$6289 N$6290 VDD VDD p L=2u W=6u
        MN186 N$6490 N$6289 GND GND n L=2u W=6u
        MP186 N$6490 N$6289 VDD VDD p L=2u W=6u
        MP193 N$6285 N$6286 N$6287 VDD p L=2u W=3u
        MP192 N$6287 N$6286 VDD VDD p L=2u W=3u
        MP191 N$6287 N$6542 VDD VDD p L=2u W=3u
        MN190 N$6299 N$6548 GND GND n L=2u W=5u
        MP185 N$6290 CK N$6490 VDD p L=2u W=6u
        MP190 GND N$6683 N$6299 VDD p L=2u W=5u
        MN189 N$6299 N$6683 N$6542 GND n L=2u W=5u
        MP77 N$1755 N$1734 VDD VDD p L=2u W=3u
        MP76 N$1752 N$1750 VDD VDD p L=2u W=3u
        MN76 N$1750 N$6255 N$1754 GND n L=2u W=3u
        MP195 N$6284 N$6542 N$6285 VDD p L=2u W=3u
        MP194 N$6284 C0 N$6287 VDD p L=2u W=3u
        MP200 N$6280 N$6542 N$6281 VDD p L=2u W=3u
        MP199 N$6281 N$6286 VDD VDD p L=2u W=3u
        MP16 N$1270 GND VDD VDD p L=2u W=3u
        MN34 N$1697 N$6233 N$1701 GND n L=2u W=3u
        MN196 N$6284 N$6542 N$6282 GND n L=2u W=3u
        MN508 N$6865 N$6777 GND GND n L=2u W=3u
        MP512 N$6777 N$6922 N$6776 VDD p L=2u W=3u
        MP511 N$6777 N$6764 N$6775 VDD p L=2u W=3u
        MP510 N$6776 N$6887 N$6775 VDD p L=2u W=3u
        MP509 N$6775 N$6887 VDD VDD p L=2u W=3u
        MP508 N$6775 N$6922 VDD VDD p L=2u W=3u
        MN510 N$6777 N$6764 N$6779 GND n L=2u W=3u
        MN474 OUT1 N$6770 GND GND n L=2u W=3u
        MP474 OUT1 N$6770 VDD VDD p L=2u W=3u
        MN405 N$6770 N$6749 N$6772 GND n L=2u W=3u
        MN404 N$6770 N$6762 N$6771 GND n L=2u W=3u
        MN403 N$6773 N$6696 GND GND n L=2u W=3u
        MN402 N$6772 N$6921 N$6773 GND n L=2u W=3u
        MN401 N$6771 N$6749 GND GND n L=2u W=3u
        MN400 N$6771 N$6696 GND GND n L=2u W=3u
        MN399 N$6771 N$6921 GND GND n L=2u W=3u
        MP405 N$6770 N$6762 N$6767 VDD p L=2u W=3u
        MP117 A2 N$6692 N$6662 VDD p L=2u W=5u
        MP338 N$6204 N$6933 N$6248 VDD p L=2u W=5u
        MN337 N$6248 N$6933 N$6921 GND n L=2u W=5u
        MP337 N$6921 N$8380 N$6248 VDD p L=2u W=5u
        MP400 N$6767 N$6921 VDD VDD p L=2u W=3u
        MP399 N$6767 N$6749 VDD VDD p L=2u W=3u
        MP398 N$6764 N$6762 VDD VDD p L=2u W=3u
        MN398 N$6762 N$6921 N$6766 GND n L=2u W=3u
        MN341 N$6252 N$6933 N$6923 GND n L=2u W=5u
        MP341 N$6923 N$8380 N$6252 VDD p L=2u W=5u
        MN340 N$6250 N$8380 N$6197 GND n L=2u W=5u
        MN509 N$6779 N$6922 GND GND n L=2u W=3u


*.ends mynand3

* Auxiliary circuit for power analysis
Cp Pav 0 100p
Rp Pav 0 100k
Fp 0 Pav Vtstp 0.003125
*Output load capacitance if you have any

*Cload1 out GND 200fF
.MODEL n NMOS LEVEL = 3
+ TOX = 200E-10 NSUB = 1E17 GAMMA = 0.5
+ PHI = 0.7 VTO = 0.8 DELTA = 3.0
+ UO = 650 ETA = 3.0E-6 THETA = 0.1
+ KP = 120E-6 VMAX = 1E5 KAPPA = 0.3
+ RSH = 0 NFS = 1E12 TPG = 1
+ XJ = 500E-9 LD = 100E-9
+ CGDO = 200E-12 CGSO = 200E-12 CGBO = 1E-10
+ CJ = 400E-6 PB = 1 MJ = 0.5
+ CJSW = 300E-12 MJSW = 0.5

.MODEL p PMOS LEVEL = 3
+ TOX = 200E-10 NSUB = 1E17 GAMMA = 0.6
+ PHI = 0.7 VTO = -0.9 DELTA = 0.1
+ UO = 250 ETA = 0 THETA = 0.1
+ KP = 40E-6 VMAX = 5E4 KAPPA = 1
+ RSH = 0 NFS = 1E12 TPG = -1
+ XJ = 500E-9 LD = 100E-9
+ CGDO = 200E-12 CGSO = 200E-12 CGBO = 1E-10
+ CJ = 400E-6 PB = 1 MJ = 0.5
+ CJSW = 300E-12 MJSW = 0.5

*Define power rails
Vddt top 0 5
Vtstp top Vdd 0
Vss GND 0 0

* Define input voltages of A and B

Vck CK 0 PWL(0 5 20N 5 20.1N 0 40N 0 40.1N 5 60N 5 60.1N 0 80N 0 80.1N 5
+ 100N 5 100.1N 0 120N 0 120.1N 5 140N 5 140.1N 0 160N 0 160.1N 5 180N 5 180.1N 0 200N 0)
Va5 A5 0 PWL(0 5 20N 5 20.1N 5 40N 5 40.1N 5 60N 5 60.1N 5 80N 5 80.1N 5
+ 100N 5 100.1N 5 120N 5 120.1N 5 140N 5 140.1N 5 160N 5 160.1N 5 180N 5 180.1N 5 200N 5)
Va0 A0 0 PWL(0 5 20N 5 20.1N 5 40N 5 40.1N 5 60N 5 60.1N 5 80N 5 80.1N 5
+ 100N 5 100.1N 5 120N 5 120.1N 5 140N 5 140.1N 5 160N 5 160.1N 5 180N 5 180.1N 5 200N 5)
Va1 A1 0 PWL(0 0 20N 0 20.1N 0 40N 0 40.1N 0 60N 0 60.1N 0 80N 0 80.1N 0
+ 100N 0 100.1N 0 120N 0 120.1N 0 140N 0 140.1N 0 160N 0 160.1N 0 180N 0 180.1N 0 200N 0)
Va2 A2 0 PWL(0 5 20N 5 20.1N 5 40N 5 40.1N 5 60N 5 60.1N 5 80N 5 80.1N 5
+ 100N 5 100.1N 5 120N 5 120.1N 5 140N 5 140.1N 5 160N 5 160.1N 5 180N 5 180.1N 5 200N 5)
Va3 A3 0 PWL(0 0 20N 0 20.1N 0 40N 0 40.1N 0 60N 0 60.1N 0 80N 0 80.1N 0
+ 100N 0 100.1N 0 120N 0 120.1N 0 140N 0 140.1N 0 160N 0 160.1N 0 180N 0 180.1N 0 200N 0)
Vrst RST 0 PWL(0 5 20N 5 20.1N 5 40N 5 40.1N 0 60N 0 60.1N 0 80N 0 80.1N 0
+ 100N 0 100.1N 0 120N 0 120.1N 0 140N 0 140.1N 0 160N 0 160.1N 0 180N 0 180.1N 0 200N 0)
Vh0 H0 0 PWL(0 5 20N 5 20.1N 5 40N 5 40.1N 5 60N 5 60.1N 5 80N 5 80.1N 5
+ 100N 5 100.1N 5 120N 5 120.1N 5 140N 5 140.1N 5 160N 5 160.1N 5 180N 5 180.1N 5 200N 5)
Vh1 H1 0 PWL(0 0 20N 0 20.1N 0 40N 0 40.1N 0 60N 0 60.1N 0 80N 0 80.1N 0
+ 100N 0 100.1N 0 120N 0 120.1N 0 140N 0 140.1N 0 160N 0 160.1N 0 180N 0 180.1N 0 200N 0)
Vh2 H2 0 PWL(0 5 20N 5 20.1N 5 40N 5 40.1N 5 60N 5 60.1N 5 80N 5 80.1N 5
+ 100N 5 100.1N 5 120N 5 120.1N 5 140N 5 140.1N 5 160N 5 160.1N 5 180N 5 180.1N 5 200N 5)
Vh3 H3 0 PWL(0 0 20N 0 20.1N 0 40N 0 40.1N 0 60N 0 60.1N 0 80N 0 80.1N 0
+ 100N 0 100.1N 0 120N 0 120.1N 0 140N 0 140.1N 0 160N 0 160.1N 0 180N 0 180.1N 0 200N 0)
Vc0 C0 0 PWL(0 0 20N 0 20.1N 0 40N 0 40.1N 0 60N 0 60.1N 0 80N 0 80.1N 0
+ 100N 0 100.1N 0 120N 0 120.1N 0 140N 0 140.1N 0 160N 0 160.1N 0 180N 0 180.1N 0 200N 0)



*Define transient simulation and probe voltage/current signals
.TRAN 20N 200N
.PROBE V(*) I(*)
.end