*
* .CONNECT statements
*
.CONNECT GND 0


* ELDO netlist generated with ICnet by 'mentor' on Fri Mar 14 2008 at 13:36:14

*
* Globals.
*
.global GND VDD

*
* MAIN CELL: Component pathname : /home/mentor/NAND/nand
*
        MN2 N$6 B GND GND n L=2u W=6u
        MN1 OUT A N$6 GND n L=2u W=6u
        MP2 OUT B VDD VDD p L=2u W=6u
        MP1 OUT A VDD VDD p L=2u W=6u
*
.end
